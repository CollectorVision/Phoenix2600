-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80db",
     9 => x"d8080b0b",
    10 => x"80dbdc08",
    11 => x"0b0b80db",
    12 => x"e0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"dbe00c0b",
    16 => x"0b80dbdc",
    17 => x"0c0b0b80",
    18 => x"dbd80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d4c0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80dbd870",
    57 => x"80e79827",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a7c9",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80db",
    65 => x"e80c9f0b",
    66 => x"80dbec0c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"dbec08ff",
    70 => x"0580dbec",
    71 => x"0c80dbec",
    72 => x"088025e8",
    73 => x"3880dbe8",
    74 => x"08ff0580",
    75 => x"dbe80c80",
    76 => x"dbe80880",
    77 => x"25d03880",
    78 => x"0b80dbec",
    79 => x"0c800b80",
    80 => x"dbe80c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80dbe808",
   100 => x"25913882",
   101 => x"c82d80db",
   102 => x"e808ff05",
   103 => x"80dbe80c",
   104 => x"838a0480",
   105 => x"dbe80880",
   106 => x"dbec0853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80dbe808",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"dbec0881",
   116 => x"0580dbec",
   117 => x"0c80dbec",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80dbec",
   121 => x"0c80dbe8",
   122 => x"08810580",
   123 => x"dbe80c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480db",
   128 => x"ec088105",
   129 => x"80dbec0c",
   130 => x"80dbec08",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80dbec",
   134 => x"0c80dbe8",
   135 => x"08810580",
   136 => x"dbe80c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"dbf00cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"dbf00c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280db",
   177 => x"f0088407",
   178 => x"80dbf00c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80d7",
   183 => x"e40c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80dbf0",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80db",
   208 => x"d80c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02f8050d",
  1093 => x"80da9408",
  1094 => x"862a7083",
  1095 => x"068207e0",
  1096 => x"0c528051",
  1097 => x"86da2d86",
  1098 => x"c72d0288",
  1099 => x"050d0402",
  1100 => x"f8050d02",
  1101 => x"8f0580f5",
  1102 => x"2d80d7ec",
  1103 => x"08525270",
  1104 => x"80dd8527",
  1105 => x"9a387171",
  1106 => x"81b72d80",
  1107 => x"d7ec0881",
  1108 => x"0580d7ec",
  1109 => x"0c80d7ec",
  1110 => x"08518071",
  1111 => x"81b72d02",
  1112 => x"88050d04",
  1113 => x"02f4050d",
  1114 => x"7470842a",
  1115 => x"708f0680",
  1116 => x"d7e80805",
  1117 => x"7080f52d",
  1118 => x"54515353",
  1119 => x"a2af2d72",
  1120 => x"8f0680d7",
  1121 => x"e8080570",
  1122 => x"80f52d52",
  1123 => x"53a2af2d",
  1124 => x"028c050d",
  1125 => x"0402f405",
  1126 => x"0d747654",
  1127 => x"52727081",
  1128 => x"055480f5",
  1129 => x"2d517072",
  1130 => x"70810554",
  1131 => x"81b72d70",
  1132 => x"ec387072",
  1133 => x"81b72d02",
  1134 => x"8c050d04",
  1135 => x"02c4050d",
  1136 => x"800b80da",
  1137 => x"9408a006",
  1138 => x"71725a40",
  1139 => x"405b810b",
  1140 => x"ec0c840b",
  1141 => x"ec0c6052",
  1142 => x"80dbf451",
  1143 => x"80cb8d2d",
  1144 => x"80dbd808",
  1145 => x"7b2e8281",
  1146 => x"3880dbf8",
  1147 => x"087bff12",
  1148 => x"575e5674",
  1149 => x"7b2e8b38",
  1150 => x"811d7581",
  1151 => x"2a565d74",
  1152 => x"f738f71d",
  1153 => x"5d815b80",
  1154 => x"762581dd",
  1155 => x"387c5274",
  1156 => x"5184a82d",
  1157 => x"80ddd052",
  1158 => x"80dbf451",
  1159 => x"80cde12d",
  1160 => x"80dbd808",
  1161 => x"802e81a7",
  1162 => x"3880ddd0",
  1163 => x"5c83ff58",
  1164 => x"7e9c387b",
  1165 => x"7081055d",
  1166 => x"80f52d77",
  1167 => x"811959e4",
  1168 => x"0ce80cff",
  1169 => x"18587780",
  1170 => x"25e938a5",
  1171 => x"d7047b70",
  1172 => x"81055d80",
  1173 => x"f52d7781",
  1174 => x"1959e40c",
  1175 => x"f4800870",
  1176 => x"72327009",
  1177 => x"81057072",
  1178 => x"079f2a51",
  1179 => x"56565b59",
  1180 => x"7d80d038",
  1181 => x"81707406",
  1182 => x"54547280",
  1183 => x"2e80c438",
  1184 => x"7380dcc8",
  1185 => x"0b80d7ec",
  1186 => x"0c80d5fc",
  1187 => x"5380dcc4",
  1188 => x"525ea395",
  1189 => x"2dff1770",
  1190 => x"5253a2e4",
  1191 => x"2d72882c",
  1192 => x"51a2e42d",
  1193 => x"a051a2af",
  1194 => x"2d7851a2",
  1195 => x"e42da051",
  1196 => x"a2af2d79",
  1197 => x"51a2e42d",
  1198 => x"80dcc452",
  1199 => x"80dc8051",
  1200 => x"a3952dff",
  1201 => x"18587780",
  1202 => x"25ff8338",
  1203 => x"a5d70480",
  1204 => x"dbd8085b",
  1205 => x"84805680",
  1206 => x"dbf45180",
  1207 => x"cdb02dfc",
  1208 => x"80168116",
  1209 => x"5656a487",
  1210 => x"0480dbf8",
  1211 => x"08f80c7d",
  1212 => x"80c23880",
  1213 => x"d6845280",
  1214 => x"dcc451a3",
  1215 => x"952d80dc",
  1216 => x"c70b80d7",
  1217 => x"ec0c7688",
  1218 => x"2c51a2e4",
  1219 => x"2d7651a2",
  1220 => x"e42da051",
  1221 => x"a2af2d80",
  1222 => x"dbf80888",
  1223 => x"2a51a2e4",
  1224 => x"2d80dbf8",
  1225 => x"0851a2e4",
  1226 => x"2d80dcc4",
  1227 => x"5280dc80",
  1228 => x"51a3952d",
  1229 => x"805186da",
  1230 => x"2d7a802e",
  1231 => x"883880d7",
  1232 => x"f051a6c9",
  1233 => x"0480d9a4",
  1234 => x"51afbc2d",
  1235 => x"7a80dbd8",
  1236 => x"0c02bc05",
  1237 => x"0d0402ec",
  1238 => x"050d80dc",
  1239 => x"c40b80d7",
  1240 => x"ec0c80dc",
  1241 => x"c4558075",
  1242 => x"81b72d80",
  1243 => x"d9c80851",
  1244 => x"a2e42dba",
  1245 => x"51a2af2d",
  1246 => x"ffb40870",
  1247 => x"982a5254",
  1248 => x"a2e42d73",
  1249 => x"902a7081",
  1250 => x"ff065253",
  1251 => x"a2e42d73",
  1252 => x"882a7081",
  1253 => x"ff065253",
  1254 => x"a2e42d73",
  1255 => x"81ff0651",
  1256 => x"a2e42d74",
  1257 => x"5280dc80",
  1258 => x"51a3952d",
  1259 => x"80d7f051",
  1260 => x"afbc2d80",
  1261 => x"d9c80884",
  1262 => x"0580d9c8",
  1263 => x"0c029405",
  1264 => x"0d04800b",
  1265 => x"80d9c80c",
  1266 => x"0402ec05",
  1267 => x"0d840bec",
  1268 => x"0cacf92d",
  1269 => x"a9ae2d81",
  1270 => x"f92d8353",
  1271 => x"acdc2d81",
  1272 => x"51858d2d",
  1273 => x"ff135372",
  1274 => x"8025f138",
  1275 => x"840bec0c",
  1276 => x"80d68851",
  1277 => x"86a02d80",
  1278 => x"c1b72d80",
  1279 => x"dbd80880",
  1280 => x"2e819438",
  1281 => x"a3bc5180",
  1282 => x"d4b72d80",
  1283 => x"d6a05280",
  1284 => x"dc8051a3",
  1285 => x"952d80d7",
  1286 => x"f051afbc",
  1287 => x"2dad9b2d",
  1288 => x"a9ba2daf",
  1289 => x"cf2d80d8",
  1290 => x"840b80f5",
  1291 => x"2d80da94",
  1292 => x"08708106",
  1293 => x"55565472",
  1294 => x"802e8538",
  1295 => x"73840754",
  1296 => x"74812a70",
  1297 => x"81065153",
  1298 => x"72802e85",
  1299 => x"38738207",
  1300 => x"5474822a",
  1301 => x"70810651",
  1302 => x"5372802e",
  1303 => x"85387381",
  1304 => x"07547483",
  1305 => x"2a708106",
  1306 => x"51537280",
  1307 => x"2e853873",
  1308 => x"88075474",
  1309 => x"842a7081",
  1310 => x"06515372",
  1311 => x"802e8538",
  1312 => x"73900754",
  1313 => x"73fc0c86",
  1314 => x"5380dbd8",
  1315 => x"08833884",
  1316 => x"5372ec0c",
  1317 => x"a8a00480",
  1318 => x"0b80dbd8",
  1319 => x"0c029405",
  1320 => x"0d047198",
  1321 => x"0c04ffb0",
  1322 => x"0880dbd8",
  1323 => x"0c04810b",
  1324 => x"ffb00c04",
  1325 => x"800bffb0",
  1326 => x"0c0402f4",
  1327 => x"050daac8",
  1328 => x"0480dbd8",
  1329 => x"0881f02e",
  1330 => x"0981068a",
  1331 => x"38810b80",
  1332 => x"da8c0caa",
  1333 => x"c80480db",
  1334 => x"d80881e0",
  1335 => x"2e098106",
  1336 => x"8a38810b",
  1337 => x"80da900c",
  1338 => x"aac80480",
  1339 => x"dbd80852",
  1340 => x"80da9008",
  1341 => x"802e8938",
  1342 => x"80dbd808",
  1343 => x"81800552",
  1344 => x"71842c72",
  1345 => x"8f065353",
  1346 => x"80da8c08",
  1347 => x"802e9a38",
  1348 => x"72842980",
  1349 => x"d9cc0572",
  1350 => x"1381712b",
  1351 => x"70097308",
  1352 => x"06730c51",
  1353 => x"5353aabc",
  1354 => x"04728429",
  1355 => x"80d9cc05",
  1356 => x"72138371",
  1357 => x"2b720807",
  1358 => x"720c5353",
  1359 => x"800b80da",
  1360 => x"900c800b",
  1361 => x"80da8c0c",
  1362 => x"80dd8851",
  1363 => x"abcf2d80",
  1364 => x"dbd808ff",
  1365 => x"24feea38",
  1366 => x"800b80db",
  1367 => x"d80c028c",
  1368 => x"050d0402",
  1369 => x"f8050d80",
  1370 => x"d9cc528f",
  1371 => x"51807270",
  1372 => x"8405540c",
  1373 => x"ff115170",
  1374 => x"8025f238",
  1375 => x"0288050d",
  1376 => x"0402f005",
  1377 => x"0d7551a9",
  1378 => x"b42d7082",
  1379 => x"2cfc0680",
  1380 => x"d9cc1172",
  1381 => x"109e0671",
  1382 => x"0870722a",
  1383 => x"70830682",
  1384 => x"742b7009",
  1385 => x"7406760c",
  1386 => x"54515657",
  1387 => x"535153a9",
  1388 => x"ae2d7180",
  1389 => x"dbd80c02",
  1390 => x"90050d04",
  1391 => x"02fc050d",
  1392 => x"72518071",
  1393 => x"0c800b84",
  1394 => x"120c0284",
  1395 => x"050d0402",
  1396 => x"f0050d75",
  1397 => x"70088412",
  1398 => x"08535353",
  1399 => x"ff547171",
  1400 => x"2ea838a9",
  1401 => x"b42d8413",
  1402 => x"08708429",
  1403 => x"14881170",
  1404 => x"087081ff",
  1405 => x"06841808",
  1406 => x"81118706",
  1407 => x"841a0c53",
  1408 => x"51555151",
  1409 => x"51a9ae2d",
  1410 => x"71547380",
  1411 => x"dbd80c02",
  1412 => x"90050d04",
  1413 => x"02f8050d",
  1414 => x"a9b42de0",
  1415 => x"08708b2a",
  1416 => x"70810651",
  1417 => x"52527080",
  1418 => x"2ea13880",
  1419 => x"dd880870",
  1420 => x"842980dd",
  1421 => x"90057381",
  1422 => x"ff06710c",
  1423 => x"515180dd",
  1424 => x"88088111",
  1425 => x"870680dd",
  1426 => x"880c5180",
  1427 => x"0b80ddb0",
  1428 => x"0ca9a62d",
  1429 => x"a9ae2d02",
  1430 => x"88050d04",
  1431 => x"02fc050d",
  1432 => x"a9b42d81",
  1433 => x"0b80ddb0",
  1434 => x"0ca9ae2d",
  1435 => x"80ddb008",
  1436 => x"5170f938",
  1437 => x"0284050d",
  1438 => x"0402fc05",
  1439 => x"0d80dd88",
  1440 => x"51abbc2d",
  1441 => x"aae32dac",
  1442 => x"9451a9a2",
  1443 => x"2d028405",
  1444 => x"0d0480dd",
  1445 => x"bc0880db",
  1446 => x"d80c0402",
  1447 => x"fc050d81",
  1448 => x"0b80da98",
  1449 => x"0c815185",
  1450 => x"8d2d0284",
  1451 => x"050d0402",
  1452 => x"fc050dad",
  1453 => x"b904a9ba",
  1454 => x"2d80f651",
  1455 => x"ab812d80",
  1456 => x"dbd808f2",
  1457 => x"3880da51",
  1458 => x"ab812d80",
  1459 => x"dbd808e6",
  1460 => x"3880dbd8",
  1461 => x"0880da98",
  1462 => x"0c80dbd8",
  1463 => x"0851858d",
  1464 => x"2d028405",
  1465 => x"0d0402ec",
  1466 => x"050d7654",
  1467 => x"8052870b",
  1468 => x"881580f5",
  1469 => x"2d565374",
  1470 => x"72248338",
  1471 => x"a0537251",
  1472 => x"83842d81",
  1473 => x"128b1580",
  1474 => x"f52d5452",
  1475 => x"727225de",
  1476 => x"38029405",
  1477 => x"0d0402f0",
  1478 => x"050d80dd",
  1479 => x"bc085481",
  1480 => x"f92d800b",
  1481 => x"80ddc00c",
  1482 => x"7308802e",
  1483 => x"81893882",
  1484 => x"0b80dbec",
  1485 => x"0c80ddc0",
  1486 => x"088f0680",
  1487 => x"dbe80c73",
  1488 => x"08527183",
  1489 => x"2e963871",
  1490 => x"83268938",
  1491 => x"71812eb0",
  1492 => x"38afa004",
  1493 => x"71852ea0",
  1494 => x"38afa004",
  1495 => x"881480f5",
  1496 => x"2d841508",
  1497 => x"80d6b053",
  1498 => x"545286a0",
  1499 => x"2d718429",
  1500 => x"13700852",
  1501 => x"52afa404",
  1502 => x"7351ade6",
  1503 => x"2dafa004",
  1504 => x"80da9408",
  1505 => x"8815082c",
  1506 => x"70810651",
  1507 => x"5271802e",
  1508 => x"883880d6",
  1509 => x"b451af9d",
  1510 => x"0480d6b8",
  1511 => x"5186a02d",
  1512 => x"84140851",
  1513 => x"86a02d80",
  1514 => x"ddc00881",
  1515 => x"0580ddc0",
  1516 => x"0c8c1454",
  1517 => x"aea80402",
  1518 => x"90050d04",
  1519 => x"7180ddbc",
  1520 => x"0cae962d",
  1521 => x"80ddc008",
  1522 => x"ff0580dd",
  1523 => x"c40c0402",
  1524 => x"e8050d80",
  1525 => x"ddbc0880",
  1526 => x"ddc80857",
  1527 => x"5580f651",
  1528 => x"ab812d80",
  1529 => x"dbd80881",
  1530 => x"2a708106",
  1531 => x"51527180",
  1532 => x"2ea438af",
  1533 => x"f904a9ba",
  1534 => x"2d80f651",
  1535 => x"ab812d80",
  1536 => x"dbd808f2",
  1537 => x"3880da98",
  1538 => x"08813270",
  1539 => x"80da980c",
  1540 => x"70525285",
  1541 => x"8d2d800b",
  1542 => x"80ddb40c",
  1543 => x"800b80dd",
  1544 => x"b80c80da",
  1545 => x"9808838d",
  1546 => x"3880da51",
  1547 => x"ab812d80",
  1548 => x"dbd80880",
  1549 => x"2e8c3880",
  1550 => x"ddb40881",
  1551 => x"800780dd",
  1552 => x"b40c80d9",
  1553 => x"51ab812d",
  1554 => x"80dbd808",
  1555 => x"802e8c38",
  1556 => x"80ddb408",
  1557 => x"80c00780",
  1558 => x"ddb40c81",
  1559 => x"9451ab81",
  1560 => x"2d80dbd8",
  1561 => x"08802e8b",
  1562 => x"3880ddb4",
  1563 => x"08900780",
  1564 => x"ddb40c81",
  1565 => x"9151ab81",
  1566 => x"2d80dbd8",
  1567 => x"08802e8b",
  1568 => x"3880ddb4",
  1569 => x"08a00780",
  1570 => x"ddb40c81",
  1571 => x"f551ab81",
  1572 => x"2d80dbd8",
  1573 => x"08802e8b",
  1574 => x"3880ddb4",
  1575 => x"08810780",
  1576 => x"ddb40c81",
  1577 => x"f251ab81",
  1578 => x"2d80dbd8",
  1579 => x"08802e8b",
  1580 => x"3880ddb4",
  1581 => x"08820780",
  1582 => x"ddb40c81",
  1583 => x"eb51ab81",
  1584 => x"2d80dbd8",
  1585 => x"08802e8b",
  1586 => x"3880ddb4",
  1587 => x"08840780",
  1588 => x"ddb40c81",
  1589 => x"f451ab81",
  1590 => x"2d80dbd8",
  1591 => x"08802e8b",
  1592 => x"3880ddb4",
  1593 => x"08880780",
  1594 => x"ddb40c80",
  1595 => x"d851ab81",
  1596 => x"2d80dbd8",
  1597 => x"08802e8c",
  1598 => x"3880ddb8",
  1599 => x"08818007",
  1600 => x"80ddb80c",
  1601 => x"9251ab81",
  1602 => x"2d80dbd8",
  1603 => x"08802e8c",
  1604 => x"3880ddb8",
  1605 => x"0880c007",
  1606 => x"80ddb80c",
  1607 => x"9451ab81",
  1608 => x"2d80dbd8",
  1609 => x"08802e8b",
  1610 => x"3880ddb8",
  1611 => x"08900780",
  1612 => x"ddb80c91",
  1613 => x"51ab812d",
  1614 => x"80dbd808",
  1615 => x"802e8b38",
  1616 => x"80ddb808",
  1617 => x"a00780dd",
  1618 => x"b80c9d51",
  1619 => x"ab812d80",
  1620 => x"dbd80880",
  1621 => x"2e8b3880",
  1622 => x"ddb80881",
  1623 => x"0780ddb8",
  1624 => x"0c9b51ab",
  1625 => x"812d80db",
  1626 => x"d808802e",
  1627 => x"8b3880dd",
  1628 => x"b8088207",
  1629 => x"80ddb80c",
  1630 => x"9c51ab81",
  1631 => x"2d80dbd8",
  1632 => x"08802e8b",
  1633 => x"3880ddb8",
  1634 => x"08840780",
  1635 => x"ddb80ca3",
  1636 => x"51ab812d",
  1637 => x"80dbd808",
  1638 => x"802e8b38",
  1639 => x"80ddb808",
  1640 => x"880780dd",
  1641 => x"b80c81fd",
  1642 => x"51ab812d",
  1643 => x"81fa51ab",
  1644 => x"812db98a",
  1645 => x"0481f551",
  1646 => x"ab812d80",
  1647 => x"dbd80881",
  1648 => x"2a708106",
  1649 => x"51527180",
  1650 => x"2eb33880",
  1651 => x"ddc40852",
  1652 => x"71802e8a",
  1653 => x"38ff1280",
  1654 => x"ddc40cb3",
  1655 => x"fd0480dd",
  1656 => x"c0081080",
  1657 => x"ddc00805",
  1658 => x"70842916",
  1659 => x"51528812",
  1660 => x"08802e89",
  1661 => x"38ff5188",
  1662 => x"12085271",
  1663 => x"2d81f251",
  1664 => x"ab812d80",
  1665 => x"dbd80881",
  1666 => x"2a708106",
  1667 => x"51527180",
  1668 => x"2eb43880",
  1669 => x"ddc008ff",
  1670 => x"1180ddc4",
  1671 => x"08565353",
  1672 => x"7372258a",
  1673 => x"38811480",
  1674 => x"ddc40cb4",
  1675 => x"c6047210",
  1676 => x"13708429",
  1677 => x"16515288",
  1678 => x"1208802e",
  1679 => x"8938fe51",
  1680 => x"88120852",
  1681 => x"712d81fd",
  1682 => x"51ab812d",
  1683 => x"80dbd808",
  1684 => x"812a7081",
  1685 => x"06515271",
  1686 => x"802eb138",
  1687 => x"80ddc408",
  1688 => x"802e8a38",
  1689 => x"800b80dd",
  1690 => x"c40cb58c",
  1691 => x"0480ddc0",
  1692 => x"081080dd",
  1693 => x"c0080570",
  1694 => x"84291651",
  1695 => x"52881208",
  1696 => x"802e8938",
  1697 => x"fd518812",
  1698 => x"0852712d",
  1699 => x"81fa51ab",
  1700 => x"812d80db",
  1701 => x"d808812a",
  1702 => x"70810651",
  1703 => x"5271802e",
  1704 => x"b13880dd",
  1705 => x"c008ff11",
  1706 => x"545280dd",
  1707 => x"c4087325",
  1708 => x"89387280",
  1709 => x"ddc40cb5",
  1710 => x"d2047110",
  1711 => x"12708429",
  1712 => x"16515288",
  1713 => x"1208802e",
  1714 => x"8938fc51",
  1715 => x"88120852",
  1716 => x"712d80dd",
  1717 => x"c4087053",
  1718 => x"5473802e",
  1719 => x"8a388c15",
  1720 => x"ff155555",
  1721 => x"b5d90482",
  1722 => x"0b80dbec",
  1723 => x"0c718f06",
  1724 => x"80dbe80c",
  1725 => x"81eb51ab",
  1726 => x"812d80db",
  1727 => x"d808812a",
  1728 => x"70810651",
  1729 => x"5271802e",
  1730 => x"ad387408",
  1731 => x"852e0981",
  1732 => x"06a43888",
  1733 => x"1580f52d",
  1734 => x"ff055271",
  1735 => x"881681b7",
  1736 => x"2d71982b",
  1737 => x"52718025",
  1738 => x"8838800b",
  1739 => x"881681b7",
  1740 => x"2d7451ad",
  1741 => x"e62d81f4",
  1742 => x"51ab812d",
  1743 => x"80dbd808",
  1744 => x"812a7081",
  1745 => x"06515271",
  1746 => x"802eb338",
  1747 => x"7408852e",
  1748 => x"098106aa",
  1749 => x"38881580",
  1750 => x"f52d8105",
  1751 => x"52718816",
  1752 => x"81b72d71",
  1753 => x"81ff068b",
  1754 => x"1680f52d",
  1755 => x"54527272",
  1756 => x"27873872",
  1757 => x"881681b7",
  1758 => x"2d7451ad",
  1759 => x"e62d80da",
  1760 => x"51ab812d",
  1761 => x"80dbd808",
  1762 => x"812a7081",
  1763 => x"06515271",
  1764 => x"802e81ad",
  1765 => x"3880ddbc",
  1766 => x"0880ddc4",
  1767 => x"08555373",
  1768 => x"802e8a38",
  1769 => x"8c13ff15",
  1770 => x"5553b79f",
  1771 => x"04720852",
  1772 => x"71822ea6",
  1773 => x"38718226",
  1774 => x"89387181",
  1775 => x"2eaa38b8",
  1776 => x"c1047183",
  1777 => x"2eb43871",
  1778 => x"842e0981",
  1779 => x"0680f238",
  1780 => x"88130851",
  1781 => x"afbc2db8",
  1782 => x"c10480dd",
  1783 => x"c4085188",
  1784 => x"13085271",
  1785 => x"2db8c104",
  1786 => x"810b8814",
  1787 => x"082b80da",
  1788 => x"94083280",
  1789 => x"da940cb8",
  1790 => x"95048813",
  1791 => x"80f52d81",
  1792 => x"058b1480",
  1793 => x"f52d5354",
  1794 => x"71742483",
  1795 => x"38805473",
  1796 => x"881481b7",
  1797 => x"2dae962d",
  1798 => x"b8c10475",
  1799 => x"08802ea4",
  1800 => x"38750851",
  1801 => x"ab812d80",
  1802 => x"dbd80881",
  1803 => x"06527180",
  1804 => x"2e8c3880",
  1805 => x"ddc40851",
  1806 => x"84160852",
  1807 => x"712d8816",
  1808 => x"5675d838",
  1809 => x"8054800b",
  1810 => x"80dbec0c",
  1811 => x"738f0680",
  1812 => x"dbe80ca0",
  1813 => x"527380dd",
  1814 => x"c4082e09",
  1815 => x"81069938",
  1816 => x"80ddc008",
  1817 => x"ff057432",
  1818 => x"70098105",
  1819 => x"7072079f",
  1820 => x"2a917131",
  1821 => x"51515353",
  1822 => x"71518384",
  1823 => x"2d811454",
  1824 => x"8e7425c2",
  1825 => x"3880da98",
  1826 => x"08527180",
  1827 => x"dbd80c02",
  1828 => x"98050d04",
  1829 => x"02f4050d",
  1830 => x"d45281ff",
  1831 => x"720c7108",
  1832 => x"5381ff72",
  1833 => x"0c72882b",
  1834 => x"83fe8006",
  1835 => x"72087081",
  1836 => x"ff065152",
  1837 => x"5381ff72",
  1838 => x"0c727107",
  1839 => x"882b7208",
  1840 => x"7081ff06",
  1841 => x"51525381",
  1842 => x"ff720c72",
  1843 => x"7107882b",
  1844 => x"72087081",
  1845 => x"ff067207",
  1846 => x"80dbd80c",
  1847 => x"5253028c",
  1848 => x"050d0402",
  1849 => x"f4050d74",
  1850 => x"767181ff",
  1851 => x"06d40c53",
  1852 => x"5380ddcc",
  1853 => x"08853871",
  1854 => x"892b5271",
  1855 => x"982ad40c",
  1856 => x"71902a70",
  1857 => x"81ff06d4",
  1858 => x"0c517188",
  1859 => x"2a7081ff",
  1860 => x"06d40c51",
  1861 => x"7181ff06",
  1862 => x"d40c7290",
  1863 => x"2a7081ff",
  1864 => x"06d40c51",
  1865 => x"d4087081",
  1866 => x"ff065151",
  1867 => x"82b8bf52",
  1868 => x"7081ff2e",
  1869 => x"09810694",
  1870 => x"3881ff0b",
  1871 => x"d40cd408",
  1872 => x"7081ff06",
  1873 => x"ff145451",
  1874 => x"5171e538",
  1875 => x"7080dbd8",
  1876 => x"0c028c05",
  1877 => x"0d0402fc",
  1878 => x"050d81c7",
  1879 => x"5181ff0b",
  1880 => x"d40cff11",
  1881 => x"51708025",
  1882 => x"f4380284",
  1883 => x"050d0402",
  1884 => x"f4050d81",
  1885 => x"ff0bd40c",
  1886 => x"93538052",
  1887 => x"87fc80c1",
  1888 => x"51b9e32d",
  1889 => x"80dbd808",
  1890 => x"8b3881ff",
  1891 => x"0bd40c81",
  1892 => x"53bb9d04",
  1893 => x"bad62dff",
  1894 => x"135372de",
  1895 => x"387280db",
  1896 => x"d80c028c",
  1897 => x"050d0402",
  1898 => x"ec050d81",
  1899 => x"0b80ddcc",
  1900 => x"0c8454d0",
  1901 => x"08708f2a",
  1902 => x"70810651",
  1903 => x"515372f3",
  1904 => x"3872d00c",
  1905 => x"bad62d80",
  1906 => x"d6bc5186",
  1907 => x"a02dd008",
  1908 => x"708f2a70",
  1909 => x"81065151",
  1910 => x"5372f338",
  1911 => x"810bd00c",
  1912 => x"b1538052",
  1913 => x"84d480c0",
  1914 => x"51b9e32d",
  1915 => x"80dbd808",
  1916 => x"812e9338",
  1917 => x"72822ebf",
  1918 => x"38ff1353",
  1919 => x"72e438ff",
  1920 => x"145473ff",
  1921 => x"ae38bad6",
  1922 => x"2d83aa52",
  1923 => x"849c80c8",
  1924 => x"51b9e32d",
  1925 => x"80dbd808",
  1926 => x"812e0981",
  1927 => x"069338b9",
  1928 => x"942d80db",
  1929 => x"d80883ff",
  1930 => x"ff065372",
  1931 => x"83aa2e9f",
  1932 => x"38baef2d",
  1933 => x"bcca0480",
  1934 => x"d6c85186",
  1935 => x"a02d8053",
  1936 => x"be9f0480",
  1937 => x"d6e05186",
  1938 => x"a02d8054",
  1939 => x"bdf00481",
  1940 => x"ff0bd40c",
  1941 => x"b154bad6",
  1942 => x"2d8fcf53",
  1943 => x"805287fc",
  1944 => x"80f751b9",
  1945 => x"e32d80db",
  1946 => x"d8085580",
  1947 => x"dbd80881",
  1948 => x"2e098106",
  1949 => x"9c3881ff",
  1950 => x"0bd40c82",
  1951 => x"0a52849c",
  1952 => x"80e951b9",
  1953 => x"e32d80db",
  1954 => x"d808802e",
  1955 => x"8d38bad6",
  1956 => x"2dff1353",
  1957 => x"72c638bd",
  1958 => x"e30481ff",
  1959 => x"0bd40c80",
  1960 => x"dbd80852",
  1961 => x"87fc80fa",
  1962 => x"51b9e32d",
  1963 => x"80dbd808",
  1964 => x"b23881ff",
  1965 => x"0bd40cd4",
  1966 => x"085381ff",
  1967 => x"0bd40c81",
  1968 => x"ff0bd40c",
  1969 => x"81ff0bd4",
  1970 => x"0c81ff0b",
  1971 => x"d40c7286",
  1972 => x"2a708106",
  1973 => x"76565153",
  1974 => x"72963880",
  1975 => x"dbd80854",
  1976 => x"bdf00473",
  1977 => x"822efedb",
  1978 => x"38ff1454",
  1979 => x"73fee738",
  1980 => x"7380ddcc",
  1981 => x"0c738b38",
  1982 => x"815287fc",
  1983 => x"80d051b9",
  1984 => x"e32d81ff",
  1985 => x"0bd40cd0",
  1986 => x"08708f2a",
  1987 => x"70810651",
  1988 => x"515372f3",
  1989 => x"3872d00c",
  1990 => x"81ff0bd4",
  1991 => x"0c815372",
  1992 => x"80dbd80c",
  1993 => x"0294050d",
  1994 => x"0402e805",
  1995 => x"0d785580",
  1996 => x"5681ff0b",
  1997 => x"d40cd008",
  1998 => x"708f2a70",
  1999 => x"81065151",
  2000 => x"5372f338",
  2001 => x"82810bd0",
  2002 => x"0c81ff0b",
  2003 => x"d40c7752",
  2004 => x"87fc80d1",
  2005 => x"51b9e32d",
  2006 => x"80dbc6df",
  2007 => x"5480dbd8",
  2008 => x"08802e8b",
  2009 => x"3880d780",
  2010 => x"5186a02d",
  2011 => x"bfc30481",
  2012 => x"ff0bd40c",
  2013 => x"d4087081",
  2014 => x"ff065153",
  2015 => x"7281fe2e",
  2016 => x"0981069e",
  2017 => x"3880ff53",
  2018 => x"b9942d80",
  2019 => x"dbd80875",
  2020 => x"70840557",
  2021 => x"0cff1353",
  2022 => x"728025ec",
  2023 => x"388156bf",
  2024 => x"a804ff14",
  2025 => x"5473c838",
  2026 => x"81ff0bd4",
  2027 => x"0c81ff0b",
  2028 => x"d40cd008",
  2029 => x"708f2a70",
  2030 => x"81065151",
  2031 => x"5372f338",
  2032 => x"72d00c75",
  2033 => x"80dbd80c",
  2034 => x"0298050d",
  2035 => x"0402e805",
  2036 => x"0d77797b",
  2037 => x"58555580",
  2038 => x"53727625",
  2039 => x"a4387470",
  2040 => x"81055680",
  2041 => x"f52d7470",
  2042 => x"81055680",
  2043 => x"f52d5252",
  2044 => x"71712e87",
  2045 => x"38815180",
  2046 => x"c0830481",
  2047 => x"1353bfd9",
  2048 => x"04805170",
  2049 => x"80dbd80c",
  2050 => x"0298050d",
  2051 => x"0402ec05",
  2052 => x"0d765574",
  2053 => x"802e80c4",
  2054 => x"389a1580",
  2055 => x"e02d5180",
  2056 => x"cebb2d80",
  2057 => x"dbd80880",
  2058 => x"dbd80880",
  2059 => x"e4800c80",
  2060 => x"dbd80854",
  2061 => x"5480e3dc",
  2062 => x"08802e9b",
  2063 => x"38941580",
  2064 => x"e02d5180",
  2065 => x"cebb2d80",
  2066 => x"dbd80890",
  2067 => x"2b83fff0",
  2068 => x"0a067075",
  2069 => x"07515372",
  2070 => x"80e4800c",
  2071 => x"80e48008",
  2072 => x"5372802e",
  2073 => x"9e3880e3",
  2074 => x"d408fe14",
  2075 => x"712980e3",
  2076 => x"e8080580",
  2077 => x"e4840c70",
  2078 => x"842b80e3",
  2079 => x"e00c5480",
  2080 => x"c1b20480",
  2081 => x"e3ec0880",
  2082 => x"e4800c80",
  2083 => x"e3f00880",
  2084 => x"e4840c80",
  2085 => x"e3dc0880",
  2086 => x"2e8c3880",
  2087 => x"e3d40884",
  2088 => x"2b5380c1",
  2089 => x"ad0480e3",
  2090 => x"f408842b",
  2091 => x"537280e3",
  2092 => x"e00c0294",
  2093 => x"050d0402",
  2094 => x"d8050d80",
  2095 => x"0b80e3dc",
  2096 => x"0c8454bb",
  2097 => x"a72d80db",
  2098 => x"d808802e",
  2099 => x"983880dd",
  2100 => x"d0528051",
  2101 => x"bea92d80",
  2102 => x"dbd80880",
  2103 => x"2e8738fe",
  2104 => x"5480c1ed",
  2105 => x"04ff1454",
  2106 => x"738024d7",
  2107 => x"38738e38",
  2108 => x"80d79051",
  2109 => x"86a02d73",
  2110 => x"5580c7cb",
  2111 => x"04805681",
  2112 => x"0b80e488",
  2113 => x"0c885380",
  2114 => x"d7a45280",
  2115 => x"de8651bf",
  2116 => x"cd2d80db",
  2117 => x"d808762e",
  2118 => x"09810689",
  2119 => x"3880dbd8",
  2120 => x"0880e488",
  2121 => x"0c885380",
  2122 => x"d7b05280",
  2123 => x"dea251bf",
  2124 => x"cd2d80db",
  2125 => x"d8088938",
  2126 => x"80dbd808",
  2127 => x"80e4880c",
  2128 => x"80e48808",
  2129 => x"802e8184",
  2130 => x"3880e196",
  2131 => x"0b80f52d",
  2132 => x"80e1970b",
  2133 => x"80f52d71",
  2134 => x"982b7190",
  2135 => x"2b0780e1",
  2136 => x"980b80f5",
  2137 => x"2d70882b",
  2138 => x"720780e1",
  2139 => x"990b80f5",
  2140 => x"2d710780",
  2141 => x"e1ce0b80",
  2142 => x"f52d80e1",
  2143 => x"cf0b80f5",
  2144 => x"2d71882b",
  2145 => x"07535f54",
  2146 => x"525a5657",
  2147 => x"557381ab",
  2148 => x"aa2e0981",
  2149 => x"06903875",
  2150 => x"5180ce8a",
  2151 => x"2d80dbd8",
  2152 => x"085680c3",
  2153 => x"b5047382",
  2154 => x"d4d52e89",
  2155 => x"3880d7bc",
  2156 => x"5180c482",
  2157 => x"0480ddd0",
  2158 => x"527551be",
  2159 => x"a92d80db",
  2160 => x"d8085580",
  2161 => x"dbd80880",
  2162 => x"2e848038",
  2163 => x"885380d7",
  2164 => x"b05280de",
  2165 => x"a251bfcd",
  2166 => x"2d80dbd8",
  2167 => x"088b3881",
  2168 => x"0b80e3dc",
  2169 => x"0c80c489",
  2170 => x"04885380",
  2171 => x"d7a45280",
  2172 => x"de8651bf",
  2173 => x"cd2d80db",
  2174 => x"d808802e",
  2175 => x"8c3880d7",
  2176 => x"d05186a0",
  2177 => x"2d80c4e8",
  2178 => x"0480e1ce",
  2179 => x"0b80f52d",
  2180 => x"547380d5",
  2181 => x"2e098106",
  2182 => x"80ce3880",
  2183 => x"e1cf0b80",
  2184 => x"f52d5473",
  2185 => x"81aa2e09",
  2186 => x"8106bd38",
  2187 => x"800b80dd",
  2188 => x"d00b80f5",
  2189 => x"2d565474",
  2190 => x"81e92e83",
  2191 => x"38815474",
  2192 => x"81eb2e8c",
  2193 => x"38805573",
  2194 => x"752e0981",
  2195 => x"0682fc38",
  2196 => x"80dddb0b",
  2197 => x"80f52d55",
  2198 => x"748e3880",
  2199 => x"dddc0b80",
  2200 => x"f52d5473",
  2201 => x"822e8738",
  2202 => x"805580c7",
  2203 => x"cb0480dd",
  2204 => x"dd0b80f5",
  2205 => x"2d7080e3",
  2206 => x"d40cff05",
  2207 => x"80e3d80c",
  2208 => x"80ddde0b",
  2209 => x"80f52d80",
  2210 => x"dddf0b80",
  2211 => x"f52d5876",
  2212 => x"05778280",
  2213 => x"29057080",
  2214 => x"e3e40c80",
  2215 => x"dde00b80",
  2216 => x"f52d7080",
  2217 => x"e3f80c80",
  2218 => x"e3dc0859",
  2219 => x"57587680",
  2220 => x"2e81b838",
  2221 => x"885380d7",
  2222 => x"b05280de",
  2223 => x"a251bfcd",
  2224 => x"2d80dbd8",
  2225 => x"08828438",
  2226 => x"80e3d408",
  2227 => x"70842b80",
  2228 => x"e3e00c70",
  2229 => x"80e3f40c",
  2230 => x"80ddf50b",
  2231 => x"80f52d80",
  2232 => x"ddf40b80",
  2233 => x"f52d7182",
  2234 => x"80290580",
  2235 => x"ddf60b80",
  2236 => x"f52d7084",
  2237 => x"80802912",
  2238 => x"80ddf70b",
  2239 => x"80f52d70",
  2240 => x"81800a29",
  2241 => x"127080e3",
  2242 => x"fc0c80e3",
  2243 => x"f8087129",
  2244 => x"80e3e408",
  2245 => x"057080e3",
  2246 => x"e80c80dd",
  2247 => x"fd0b80f5",
  2248 => x"2d80ddfc",
  2249 => x"0b80f52d",
  2250 => x"71828029",
  2251 => x"0580ddfe",
  2252 => x"0b80f52d",
  2253 => x"70848080",
  2254 => x"291280dd",
  2255 => x"ff0b80f5",
  2256 => x"2d70982b",
  2257 => x"81f00a06",
  2258 => x"72057080",
  2259 => x"e3ec0cfe",
  2260 => x"117e2977",
  2261 => x"0580e3f0",
  2262 => x"0c525952",
  2263 => x"43545e51",
  2264 => x"5259525d",
  2265 => x"57595780",
  2266 => x"c7c30480",
  2267 => x"dde20b80",
  2268 => x"f52d80dd",
  2269 => x"e10b80f5",
  2270 => x"2d718280",
  2271 => x"29057080",
  2272 => x"e3e00c70",
  2273 => x"a02983ff",
  2274 => x"0570892a",
  2275 => x"7080e3f4",
  2276 => x"0c80dde7",
  2277 => x"0b80f52d",
  2278 => x"80dde60b",
  2279 => x"80f52d71",
  2280 => x"82802905",
  2281 => x"7080e3fc",
  2282 => x"0c7b7129",
  2283 => x"1e7080e3",
  2284 => x"f00c7d80",
  2285 => x"e3ec0c73",
  2286 => x"0580e3e8",
  2287 => x"0c555e51",
  2288 => x"51555580",
  2289 => x"5180c08d",
  2290 => x"2d815574",
  2291 => x"80dbd80c",
  2292 => x"02a8050d",
  2293 => x"0402ec05",
  2294 => x"0d767087",
  2295 => x"2c7180ff",
  2296 => x"06555654",
  2297 => x"80e3dc08",
  2298 => x"8a387388",
  2299 => x"2c7481ff",
  2300 => x"06545580",
  2301 => x"ddd05280",
  2302 => x"e3e40815",
  2303 => x"51bea92d",
  2304 => x"80dbd808",
  2305 => x"5480dbd8",
  2306 => x"08802ebb",
  2307 => x"3880e3dc",
  2308 => x"08802e9c",
  2309 => x"38728429",
  2310 => x"80ddd005",
  2311 => x"70085253",
  2312 => x"80ce8a2d",
  2313 => x"80dbd808",
  2314 => x"f00a0653",
  2315 => x"80c8c504",
  2316 => x"721080dd",
  2317 => x"d0057080",
  2318 => x"e02d5253",
  2319 => x"80cebb2d",
  2320 => x"80dbd808",
  2321 => x"53725473",
  2322 => x"80dbd80c",
  2323 => x"0294050d",
  2324 => x"0402e005",
  2325 => x"0d797084",
  2326 => x"2c80e484",
  2327 => x"0805718f",
  2328 => x"06525553",
  2329 => x"728a3880",
  2330 => x"ddd05273",
  2331 => x"51bea92d",
  2332 => x"72a02980",
  2333 => x"ddd00554",
  2334 => x"807480f5",
  2335 => x"2d565374",
  2336 => x"732e8338",
  2337 => x"81537481",
  2338 => x"e52e81f5",
  2339 => x"38817074",
  2340 => x"06545872",
  2341 => x"802e81e9",
  2342 => x"388b1480",
  2343 => x"f52d7083",
  2344 => x"2a790658",
  2345 => x"56769c38",
  2346 => x"80da9c08",
  2347 => x"53728938",
  2348 => x"7280e1d0",
  2349 => x"0b81b72d",
  2350 => x"7680da9c",
  2351 => x"0c735380",
  2352 => x"cb830475",
  2353 => x"8f2e0981",
  2354 => x"0681b638",
  2355 => x"749f068d",
  2356 => x"2980e1c3",
  2357 => x"11515381",
  2358 => x"1480f52d",
  2359 => x"73708105",
  2360 => x"5581b72d",
  2361 => x"831480f5",
  2362 => x"2d737081",
  2363 => x"055581b7",
  2364 => x"2d851480",
  2365 => x"f52d7370",
  2366 => x"81055581",
  2367 => x"b72d8714",
  2368 => x"80f52d73",
  2369 => x"70810555",
  2370 => x"81b72d89",
  2371 => x"1480f52d",
  2372 => x"73708105",
  2373 => x"5581b72d",
  2374 => x"8e1480f5",
  2375 => x"2d737081",
  2376 => x"055581b7",
  2377 => x"2d901480",
  2378 => x"f52d7370",
  2379 => x"81055581",
  2380 => x"b72d9214",
  2381 => x"80f52d73",
  2382 => x"70810555",
  2383 => x"81b72d94",
  2384 => x"1480f52d",
  2385 => x"73708105",
  2386 => x"5581b72d",
  2387 => x"961480f5",
  2388 => x"2d737081",
  2389 => x"055581b7",
  2390 => x"2d981480",
  2391 => x"f52d7370",
  2392 => x"81055581",
  2393 => x"b72d9c14",
  2394 => x"80f52d73",
  2395 => x"70810555",
  2396 => x"81b72d9e",
  2397 => x"1480f52d",
  2398 => x"7381b72d",
  2399 => x"7780da9c",
  2400 => x"0c805372",
  2401 => x"80dbd80c",
  2402 => x"02a0050d",
  2403 => x"0402cc05",
  2404 => x"0d7e605e",
  2405 => x"5a800b80",
  2406 => x"e4800880",
  2407 => x"e4840859",
  2408 => x"5c568058",
  2409 => x"80e3e008",
  2410 => x"782e81bc",
  2411 => x"38778f06",
  2412 => x"a0175754",
  2413 => x"73913880",
  2414 => x"ddd05276",
  2415 => x"51811757",
  2416 => x"bea92d80",
  2417 => x"ddd05680",
  2418 => x"7680f52d",
  2419 => x"56547474",
  2420 => x"2e833881",
  2421 => x"547481e5",
  2422 => x"2e818138",
  2423 => x"81707506",
  2424 => x"555c7380",
  2425 => x"2e80f538",
  2426 => x"8b1680f5",
  2427 => x"2d980659",
  2428 => x"7880e938",
  2429 => x"8b537c52",
  2430 => x"7551bfcd",
  2431 => x"2d80dbd8",
  2432 => x"0880d938",
  2433 => x"9c160851",
  2434 => x"80ce8a2d",
  2435 => x"80dbd808",
  2436 => x"841b0c9a",
  2437 => x"1680e02d",
  2438 => x"5180cebb",
  2439 => x"2d80dbd8",
  2440 => x"0880dbd8",
  2441 => x"08881c0c",
  2442 => x"80dbd808",
  2443 => x"555580e3",
  2444 => x"dc08802e",
  2445 => x"9a389416",
  2446 => x"80e02d51",
  2447 => x"80cebb2d",
  2448 => x"80dbd808",
  2449 => x"902b83ff",
  2450 => x"f00a0670",
  2451 => x"16515473",
  2452 => x"881b0c78",
  2453 => x"7a0c7b54",
  2454 => x"80cda604",
  2455 => x"81185880",
  2456 => x"e3e00878",
  2457 => x"26fec638",
  2458 => x"80e3dc08",
  2459 => x"802eb538",
  2460 => x"7a5180c7",
  2461 => x"d52d80db",
  2462 => x"d80880db",
  2463 => x"d80880ff",
  2464 => x"fffff806",
  2465 => x"555b7380",
  2466 => x"fffffff8",
  2467 => x"2e963880",
  2468 => x"dbd808fe",
  2469 => x"0580e3d4",
  2470 => x"082980e3",
  2471 => x"e8080557",
  2472 => x"80cba204",
  2473 => x"80547380",
  2474 => x"dbd80c02",
  2475 => x"b4050d04",
  2476 => x"02f4050d",
  2477 => x"74700881",
  2478 => x"05710c70",
  2479 => x"0880e3d8",
  2480 => x"08065353",
  2481 => x"71903888",
  2482 => x"13085180",
  2483 => x"c7d52d80",
  2484 => x"dbd80888",
  2485 => x"140c810b",
  2486 => x"80dbd80c",
  2487 => x"028c050d",
  2488 => x"0402f005",
  2489 => x"0d758811",
  2490 => x"08fe0580",
  2491 => x"e3d40829",
  2492 => x"80e3e808",
  2493 => x"11720880",
  2494 => x"e3d80806",
  2495 => x"05795553",
  2496 => x"5454bea9",
  2497 => x"2d029005",
  2498 => x"0d0402f4",
  2499 => x"050d7470",
  2500 => x"882a83fe",
  2501 => x"80067072",
  2502 => x"982a0772",
  2503 => x"882b87fc",
  2504 => x"80800673",
  2505 => x"982b81f0",
  2506 => x"0a067173",
  2507 => x"070780db",
  2508 => x"d80c5651",
  2509 => x"5351028c",
  2510 => x"050d0402",
  2511 => x"f8050d02",
  2512 => x"8e0580f5",
  2513 => x"2d74882b",
  2514 => x"077083ff",
  2515 => x"ff0680db",
  2516 => x"d80c5102",
  2517 => x"88050d04",
  2518 => x"02f4050d",
  2519 => x"74767853",
  2520 => x"54528071",
  2521 => x"25973872",
  2522 => x"70810554",
  2523 => x"80f52d72",
  2524 => x"70810554",
  2525 => x"81b72dff",
  2526 => x"115170eb",
  2527 => x"38807281",
  2528 => x"b72d028c",
  2529 => x"050d0402",
  2530 => x"e8050d77",
  2531 => x"56807056",
  2532 => x"54737624",
  2533 => x"b73880e3",
  2534 => x"e008742e",
  2535 => x"af387351",
  2536 => x"80c8d12d",
  2537 => x"80dbd808",
  2538 => x"80dbd808",
  2539 => x"09810570",
  2540 => x"80dbd808",
  2541 => x"079f2a77",
  2542 => x"05811757",
  2543 => x"57535374",
  2544 => x"76248938",
  2545 => x"80e3e008",
  2546 => x"7426d338",
  2547 => x"7280dbd8",
  2548 => x"0c029805",
  2549 => x"0d0402f0",
  2550 => x"050d80db",
  2551 => x"d4081651",
  2552 => x"80cf872d",
  2553 => x"80dbd808",
  2554 => x"802ea038",
  2555 => x"8b5380db",
  2556 => x"d8085280",
  2557 => x"e1d05180",
  2558 => x"ced82d80",
  2559 => x"e48c0854",
  2560 => x"73802e87",
  2561 => x"3880e1d0",
  2562 => x"51732d02",
  2563 => x"90050d04",
  2564 => x"02dc050d",
  2565 => x"80705a55",
  2566 => x"7480dbd4",
  2567 => x"0825b538",
  2568 => x"80e3e008",
  2569 => x"752ead38",
  2570 => x"785180c8",
  2571 => x"d12d80db",
  2572 => x"d8080981",
  2573 => x"057080db",
  2574 => x"d808079f",
  2575 => x"2a760581",
  2576 => x"1b5b5654",
  2577 => x"7480dbd4",
  2578 => x"08258938",
  2579 => x"80e3e008",
  2580 => x"7926d538",
  2581 => x"80557880",
  2582 => x"e3e00827",
  2583 => x"81e43878",
  2584 => x"5180c8d1",
  2585 => x"2d80dbd8",
  2586 => x"08802e81",
  2587 => x"b43880db",
  2588 => x"d8088b05",
  2589 => x"80f52d70",
  2590 => x"842a7081",
  2591 => x"06771078",
  2592 => x"842b80e1",
  2593 => x"d00b80f5",
  2594 => x"2d5c5c53",
  2595 => x"51555673",
  2596 => x"802e80ce",
  2597 => x"38741682",
  2598 => x"2b80d2e6",
  2599 => x"0b80daa8",
  2600 => x"120c5477",
  2601 => x"75311080",
  2602 => x"e4901155",
  2603 => x"56907470",
  2604 => x"81055681",
  2605 => x"b72da074",
  2606 => x"81b72d76",
  2607 => x"81ff0681",
  2608 => x"16585473",
  2609 => x"802e8b38",
  2610 => x"9c5380e1",
  2611 => x"d05280d1",
  2612 => x"d9048b53",
  2613 => x"80dbd808",
  2614 => x"5280e492",
  2615 => x"165180d2",
  2616 => x"97047416",
  2617 => x"822b80cf",
  2618 => x"d60b80da",
  2619 => x"a8120c54",
  2620 => x"7681ff06",
  2621 => x"81165854",
  2622 => x"73802e8b",
  2623 => x"389c5380",
  2624 => x"e1d05280",
  2625 => x"d28e048b",
  2626 => x"5380dbd8",
  2627 => x"08527775",
  2628 => x"311080e4",
  2629 => x"90055176",
  2630 => x"5580ced8",
  2631 => x"2d80d2b6",
  2632 => x"04749029",
  2633 => x"75317010",
  2634 => x"80e49005",
  2635 => x"515480db",
  2636 => x"d8087481",
  2637 => x"b72d8119",
  2638 => x"59748b24",
  2639 => x"a43880d0",
  2640 => x"d6047490",
  2641 => x"29753170",
  2642 => x"1080e490",
  2643 => x"058c7731",
  2644 => x"57515480",
  2645 => x"7481b72d",
  2646 => x"9e14ff16",
  2647 => x"565474f3",
  2648 => x"3802a405",
  2649 => x"0d0402fc",
  2650 => x"050d80db",
  2651 => x"d4081351",
  2652 => x"80cf872d",
  2653 => x"80dbd808",
  2654 => x"802e8a38",
  2655 => x"80dbd808",
  2656 => x"5180c08d",
  2657 => x"2d800b80",
  2658 => x"dbd40c80",
  2659 => x"d0902dae",
  2660 => x"962d0284",
  2661 => x"050d0402",
  2662 => x"fc050d72",
  2663 => x"5170fd2e",
  2664 => x"b23870fd",
  2665 => x"248b3870",
  2666 => x"fc2e80d0",
  2667 => x"3880d486",
  2668 => x"0470fe2e",
  2669 => x"b93870ff",
  2670 => x"2e098106",
  2671 => x"80c83880",
  2672 => x"dbd40851",
  2673 => x"70802ebe",
  2674 => x"38ff1180",
  2675 => x"dbd40c80",
  2676 => x"d4860480",
  2677 => x"dbd408f0",
  2678 => x"057080db",
  2679 => x"d40c5170",
  2680 => x"8025a338",
  2681 => x"800b80db",
  2682 => x"d40c80d4",
  2683 => x"860480db",
  2684 => x"d4088105",
  2685 => x"80dbd40c",
  2686 => x"80d48604",
  2687 => x"80dbd408",
  2688 => x"900580db",
  2689 => x"d40c80d0",
  2690 => x"902dae96",
  2691 => x"2d028405",
  2692 => x"0d0402fc",
  2693 => x"050d800b",
  2694 => x"80dbd40c",
  2695 => x"80d0902d",
  2696 => x"ad922d80",
  2697 => x"dbd80880",
  2698 => x"dbc40c80",
  2699 => x"daa051af",
  2700 => x"bc2d0284",
  2701 => x"050d0471",
  2702 => x"80e48c0c",
  2703 => x"04000000",
  2704 => x"00ffffff",
  2705 => x"ff00ffff",
  2706 => x"ffff00ff",
  2707 => x"ffffff00",
  2708 => x"30313233",
  2709 => x"34353637",
  2710 => x"38394142",
  2711 => x"43444546",
  2712 => x"00000000",
  2713 => x"44656275",
  2714 => x"67000000",
  2715 => x"52657365",
  2716 => x"74000000",
  2717 => x"5363616e",
  2718 => x"6c696e65",
  2719 => x"73000000",
  2720 => x"50414c20",
  2721 => x"2f204e54",
  2722 => x"53430000",
  2723 => x"436f6c6f",
  2724 => x"72000000",
  2725 => x"44696666",
  2726 => x"6963756c",
  2727 => x"74792041",
  2728 => x"00000000",
  2729 => x"44696666",
  2730 => x"6963756c",
  2731 => x"74792042",
  2732 => x"00000000",
  2733 => x"524f4d00",
  2734 => x"626f6f74",
  2735 => x"00000000",
  2736 => x"53656c65",
  2737 => x"63740000",
  2738 => x"53746172",
  2739 => x"74000000",
  2740 => x"4c6f6164",
  2741 => x"20524f4d",
  2742 => x"20100000",
  2743 => x"45786974",
  2744 => x"00000000",
  2745 => x"524f4d20",
  2746 => x"6c6f6164",
  2747 => x"696e6720",
  2748 => x"6661696c",
  2749 => x"65640000",
  2750 => x"4f4b0000",
  2751 => x"45525220",
  2752 => x"00000000",
  2753 => x"4f4b2000",
  2754 => x"496e6974",
  2755 => x"69616c69",
  2756 => x"7a696e67",
  2757 => x"20534420",
  2758 => x"63617264",
  2759 => x"0a000000",
  2760 => x"436f6c6c",
  2761 => x"6563746f",
  2762 => x"72566973",
  2763 => x"696f6e00",
  2764 => x"16200000",
  2765 => x"14200000",
  2766 => x"15200000",
  2767 => x"53442069",
  2768 => x"6e69742e",
  2769 => x"2e2e0a00",
  2770 => x"53442063",
  2771 => x"61726420",
  2772 => x"72657365",
  2773 => x"74206661",
  2774 => x"696c6564",
  2775 => x"210a0000",
  2776 => x"53444843",
  2777 => x"20657272",
  2778 => x"6f72210a",
  2779 => x"00000000",
  2780 => x"57726974",
  2781 => x"65206661",
  2782 => x"696c6564",
  2783 => x"0a000000",
  2784 => x"52656164",
  2785 => x"20666169",
  2786 => x"6c65640a",
  2787 => x"00000000",
  2788 => x"43617264",
  2789 => x"20696e69",
  2790 => x"74206661",
  2791 => x"696c6564",
  2792 => x"0a000000",
  2793 => x"46415431",
  2794 => x"36202020",
  2795 => x"00000000",
  2796 => x"46415433",
  2797 => x"32202020",
  2798 => x"00000000",
  2799 => x"4e6f2070",
  2800 => x"61727469",
  2801 => x"74696f6e",
  2802 => x"20736967",
  2803 => x"0a000000",
  2804 => x"42616420",
  2805 => x"70617274",
  2806 => x"0a000000",
  2807 => x"4261636b",
  2808 => x"00000000",
  2809 => x"00000002",
  2810 => x"00002a50",
  2811 => x"00002e44",
  2812 => x"00000002",
  2813 => x"00002e00",
  2814 => x"000013c2",
  2815 => x"00000002",
  2816 => x"00002a64",
  2817 => x"00001356",
  2818 => x"00000002",
  2819 => x"00002a6c",
  2820 => x"0000035a",
  2821 => x"00000001",
  2822 => x"00002a74",
  2823 => x"00000000",
  2824 => x"00000001",
  2825 => x"00002a80",
  2826 => x"00000001",
  2827 => x"00000001",
  2828 => x"00002a8c",
  2829 => x"00000002",
  2830 => x"00000001",
  2831 => x"00002a94",
  2832 => x"00000003",
  2833 => x"00000001",
  2834 => x"00002aa4",
  2835 => x"00000004",
  2836 => x"00000001",
  2837 => x"00002ab4",
  2838 => x"00000006",
  2839 => x"00000002",
  2840 => x"00002ab8",
  2841 => x"00001110",
  2842 => x"00000002",
  2843 => x"00002ac0",
  2844 => x"0000036e",
  2845 => x"00000002",
  2846 => x"00002ac8",
  2847 => x"00000a3f",
  2848 => x"00000002",
  2849 => x"00002ad0",
  2850 => x"00002a12",
  2851 => x"00000002",
  2852 => x"00002adc",
  2853 => x"000016af",
  2854 => x"00000000",
  2855 => x"00000000",
  2856 => x"00000000",
  2857 => x"00000004",
  2858 => x"00002ae4",
  2859 => x"00002ca4",
  2860 => x"00000004",
  2861 => x"00002af8",
  2862 => x"00002bf0",
  2863 => x"00000000",
  2864 => x"00000000",
  2865 => x"00000000",
  2866 => x"00000000",
  2867 => x"00000000",
  2868 => x"00000000",
  2869 => x"00000000",
  2870 => x"00000000",
  2871 => x"00000000",
  2872 => x"00000000",
  2873 => x"00000000",
  2874 => x"00000000",
  2875 => x"00000000",
  2876 => x"00000000",
  2877 => x"00000000",
  2878 => x"00000000",
  2879 => x"00000000",
  2880 => x"00000000",
  2881 => x"00000000",
  2882 => x"00000000",
  2883 => x"00000000",
  2884 => x"00000000",
  2885 => x"00000006",
  2886 => x"00000000",
  2887 => x"00000000",
  2888 => x"00000002",
  2889 => x"00003210",
  2890 => x"000027d6",
  2891 => x"00000002",
  2892 => x"0000322e",
  2893 => x"000027d6",
  2894 => x"00000002",
  2895 => x"0000324c",
  2896 => x"000027d6",
  2897 => x"00000002",
  2898 => x"0000326a",
  2899 => x"000027d6",
  2900 => x"00000002",
  2901 => x"00003288",
  2902 => x"000027d6",
  2903 => x"00000002",
  2904 => x"000032a6",
  2905 => x"000027d6",
  2906 => x"00000002",
  2907 => x"000032c4",
  2908 => x"000027d6",
  2909 => x"00000002",
  2910 => x"000032e2",
  2911 => x"000027d6",
  2912 => x"00000002",
  2913 => x"00003300",
  2914 => x"000027d6",
  2915 => x"00000002",
  2916 => x"0000331e",
  2917 => x"000027d6",
  2918 => x"00000002",
  2919 => x"0000333c",
  2920 => x"000027d6",
  2921 => x"00000002",
  2922 => x"0000335a",
  2923 => x"000027d6",
  2924 => x"00000002",
  2925 => x"00003378",
  2926 => x"000027d6",
  2927 => x"00000004",
  2928 => x"00002bdc",
  2929 => x"00000000",
  2930 => x"00000000",
  2931 => x"00000000",
  2932 => x"00002997",
  2933 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

