-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80dc",
     9 => x"bc080b0b",
    10 => x"80dcc008",
    11 => x"0b0b80dc",
    12 => x"c4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"dcc40c0b",
    16 => x"0b80dcc0",
    17 => x"0c0b0b80",
    18 => x"dcbc0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d4e8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80dcbc70",
    57 => x"80e7fc27",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a5ed",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80dc",
    65 => x"cc0c9f0b",
    66 => x"80dcd00c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"dcd008ff",
    70 => x"0580dcd0",
    71 => x"0c80dcd0",
    72 => x"088025e8",
    73 => x"3880dccc",
    74 => x"08ff0580",
    75 => x"dccc0c80",
    76 => x"dccc0880",
    77 => x"25d03880",
    78 => x"0b80dcd0",
    79 => x"0c800b80",
    80 => x"dccc0c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80dccc08",
   100 => x"25913882",
   101 => x"c82d80dc",
   102 => x"cc08ff05",
   103 => x"80dccc0c",
   104 => x"838a0480",
   105 => x"dccc0880",
   106 => x"dcd00853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80dccc08",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"dcd00881",
   116 => x"0580dcd0",
   117 => x"0c80dcd0",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80dcd0",
   121 => x"0c80dccc",
   122 => x"08810580",
   123 => x"dccc0c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480dc",
   128 => x"d0088105",
   129 => x"80dcd00c",
   130 => x"80dcd008",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80dcd0",
   134 => x"0c80dccc",
   135 => x"08810580",
   136 => x"dccc0c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"dcd40cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"dcd40c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280dc",
   177 => x"d4088407",
   178 => x"80dcd40c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80d8",
   183 => x"a40c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80dcd4",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80dc",
   208 => x"bc0c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02f8050d",
  1093 => x"028f0580",
  1094 => x"f52d80d8",
  1095 => x"ac085252",
  1096 => x"7080dde9",
  1097 => x"279a3871",
  1098 => x"7181b72d",
  1099 => x"80d8ac08",
  1100 => x"810580d8",
  1101 => x"ac0c80d8",
  1102 => x"ac085180",
  1103 => x"7181b72d",
  1104 => x"0288050d",
  1105 => x"0402f405",
  1106 => x"0d747084",
  1107 => x"2a708f06",
  1108 => x"80d8a808",
  1109 => x"057080f5",
  1110 => x"2d545153",
  1111 => x"53a2902d",
  1112 => x"728f0680",
  1113 => x"d8a80805",
  1114 => x"7080f52d",
  1115 => x"5253a290",
  1116 => x"2d028c05",
  1117 => x"0d0402f4",
  1118 => x"050d7476",
  1119 => x"54527270",
  1120 => x"81055480",
  1121 => x"f52d5170",
  1122 => x"72708105",
  1123 => x"5481b72d",
  1124 => x"70ec3870",
  1125 => x"7281b72d",
  1126 => x"028c050d",
  1127 => x"0402d005",
  1128 => x"0d800b80",
  1129 => x"daf80881",
  1130 => x"8006715d",
  1131 => x"5d59810b",
  1132 => x"ec0c840b",
  1133 => x"ec0c7d52",
  1134 => x"80dcd851",
  1135 => x"80cbb62d",
  1136 => x"80dcbc08",
  1137 => x"792e80ff",
  1138 => x"3880dcdc",
  1139 => x"0879ff12",
  1140 => x"57595774",
  1141 => x"792e8b38",
  1142 => x"81187581",
  1143 => x"2a565874",
  1144 => x"f738f718",
  1145 => x"58815980",
  1146 => x"772580db",
  1147 => x"38775274",
  1148 => x"5184a82d",
  1149 => x"80deb452",
  1150 => x"80dcd851",
  1151 => x"80ce8a2d",
  1152 => x"80dcbc08",
  1153 => x"802ea638",
  1154 => x"80deb45a",
  1155 => x"7ba73883",
  1156 => x"ff567970",
  1157 => x"81055b80",
  1158 => x"f52d7b81",
  1159 => x"1d5de40c",
  1160 => x"e80cff16",
  1161 => x"56758025",
  1162 => x"e938a4b5",
  1163 => x"0480dcbc",
  1164 => x"08598480",
  1165 => x"5780dcd8",
  1166 => x"5180cdd9",
  1167 => x"2dfc8017",
  1168 => x"81165657",
  1169 => x"a3e70480",
  1170 => x"dcdc08f8",
  1171 => x"0c810be0",
  1172 => x"0c805186",
  1173 => x"da2d86c7",
  1174 => x"2d78802e",
  1175 => x"883880d8",
  1176 => x"b051a4e9",
  1177 => x"0480d9f0",
  1178 => x"51afe42d",
  1179 => x"7880dcbc",
  1180 => x"0c02b005",
  1181 => x"0d0402ec",
  1182 => x"050d80dd",
  1183 => x"a80b80d8",
  1184 => x"ac0c80dd",
  1185 => x"a8538073",
  1186 => x"81b72d80",
  1187 => x"da940851",
  1188 => x"a2c52dba",
  1189 => x"51a2902d",
  1190 => x"ffb408ff",
  1191 => x"b8087098",
  1192 => x"2a535155",
  1193 => x"a2c52d74",
  1194 => x"902a7081",
  1195 => x"ff065254",
  1196 => x"a2c52d74",
  1197 => x"882a7081",
  1198 => x"ff065254",
  1199 => x"a2c52d74",
  1200 => x"81ff0651",
  1201 => x"a2c52d72",
  1202 => x"5280dce4",
  1203 => x"51a2f62d",
  1204 => x"80d8b051",
  1205 => x"afe42d80",
  1206 => x"da940884",
  1207 => x"0580da94",
  1208 => x"0c029405",
  1209 => x"0d04800b",
  1210 => x"80da940c",
  1211 => x"0402ec05",
  1212 => x"0d840bec",
  1213 => x"0cada12d",
  1214 => x"a8872d81",
  1215 => x"f92d8353",
  1216 => x"ad842d81",
  1217 => x"51858d2d",
  1218 => x"ff135372",
  1219 => x"8025f138",
  1220 => x"840bec0c",
  1221 => x"80d6c851",
  1222 => x"86a02d80",
  1223 => x"c1e02d80",
  1224 => x"dcbc0880",
  1225 => x"2e81c938",
  1226 => x"a39d5180",
  1227 => x"d4e02d80",
  1228 => x"d6e05280",
  1229 => x"dce451a2",
  1230 => x"f62d80d8",
  1231 => x"b051afe4",
  1232 => x"2dadc32d",
  1233 => x"a8d82daf",
  1234 => x"f72d80d8",
  1235 => x"c40b80f5",
  1236 => x"2d80daf8",
  1237 => x"08708106",
  1238 => x"55565472",
  1239 => x"802e8538",
  1240 => x"73840754",
  1241 => x"74812a70",
  1242 => x"81065153",
  1243 => x"72802e85",
  1244 => x"38738207",
  1245 => x"5474822a",
  1246 => x"70810651",
  1247 => x"5372802e",
  1248 => x"85387381",
  1249 => x"07547483",
  1250 => x"2a708106",
  1251 => x"51537280",
  1252 => x"2e853873",
  1253 => x"88075474",
  1254 => x"842a7081",
  1255 => x"06515372",
  1256 => x"802e8538",
  1257 => x"73900754",
  1258 => x"74852a70",
  1259 => x"81065153",
  1260 => x"72802e85",
  1261 => x"3873a007",
  1262 => x"5474882a",
  1263 => x"70810651",
  1264 => x"5372802e",
  1265 => x"86387380",
  1266 => x"c0075474",
  1267 => x"892a7081",
  1268 => x"06515372",
  1269 => x"802e8638",
  1270 => x"73818007",
  1271 => x"5473fc0c",
  1272 => x"865380dc",
  1273 => x"bc088338",
  1274 => x"845372ec",
  1275 => x"0ca6c404",
  1276 => x"800b80dc",
  1277 => x"bc0c0294",
  1278 => x"050d0471",
  1279 => x"980c04ff",
  1280 => x"b00880dc",
  1281 => x"bc0c0481",
  1282 => x"0bffb00c",
  1283 => x"04800bff",
  1284 => x"b00c0402",
  1285 => x"f8050dff",
  1286 => x"b408709f",
  1287 => x"ff065151",
  1288 => x"7080dae8",
  1289 => x"082e8c38",
  1290 => x"7080dae8",
  1291 => x"0c800b80",
  1292 => x"dae40c80",
  1293 => x"dae40851",
  1294 => x"81527087",
  1295 => x"e82e8f38",
  1296 => x"7087e824",
  1297 => x"87387111",
  1298 => x"80dae40c",
  1299 => x"80527180",
  1300 => x"dcbc0c02",
  1301 => x"88050d04",
  1302 => x"02e0050d",
  1303 => x"a9e60480",
  1304 => x"dcbc0881",
  1305 => x"f02e0981",
  1306 => x"068a3881",
  1307 => x"0b80daf0",
  1308 => x"0ca9e604",
  1309 => x"80dcbc08",
  1310 => x"81e02e09",
  1311 => x"81068a38",
  1312 => x"810b80da",
  1313 => x"f40ca9e6",
  1314 => x"0480dcbc",
  1315 => x"085280da",
  1316 => x"f408802e",
  1317 => x"893880dc",
  1318 => x"bc088180",
  1319 => x"05527184",
  1320 => x"2c728f06",
  1321 => x"535380da",
  1322 => x"f008802e",
  1323 => x"9a387284",
  1324 => x"2980da98",
  1325 => x"05721381",
  1326 => x"712b7009",
  1327 => x"73080673",
  1328 => x"0c515353",
  1329 => x"a9da0472",
  1330 => x"842980da",
  1331 => x"98057213",
  1332 => x"83712b72",
  1333 => x"0807720c",
  1334 => x"5353800b",
  1335 => x"80daf40c",
  1336 => x"800b80da",
  1337 => x"f00c80dd",
  1338 => x"ec51abf7",
  1339 => x"2d80dcbc",
  1340 => x"08ff24fe",
  1341 => x"ea38a893",
  1342 => x"2d80dcbc",
  1343 => x"08802e80",
  1344 => x"ff388156",
  1345 => x"800b80da",
  1346 => x"ec0880da",
  1347 => x"e80880da",
  1348 => x"f0085759",
  1349 => x"59557776",
  1350 => x"06777706",
  1351 => x"54527173",
  1352 => x"2e80c438",
  1353 => x"7280dad8",
  1354 => x"1680f52d",
  1355 => x"70842c71",
  1356 => x"8f065255",
  1357 => x"53547380",
  1358 => x"2e9a3872",
  1359 => x"842980da",
  1360 => x"98057213",
  1361 => x"81712b70",
  1362 => x"09730806",
  1363 => x"730c5153",
  1364 => x"53aae704",
  1365 => x"72842980",
  1366 => x"da980572",
  1367 => x"1383712b",
  1368 => x"72080772",
  1369 => x"0c535375",
  1370 => x"10811656",
  1371 => x"568b7525",
  1372 => x"ffa43873",
  1373 => x"80daf00c",
  1374 => x"80dae808",
  1375 => x"80daec0c",
  1376 => x"800b80dc",
  1377 => x"bc0c02a0",
  1378 => x"050d0402",
  1379 => x"f8050d80",
  1380 => x"da98528f",
  1381 => x"51807270",
  1382 => x"8405540c",
  1383 => x"ff115170",
  1384 => x"8025f238",
  1385 => x"0288050d",
  1386 => x"0402f005",
  1387 => x"0d7551a8",
  1388 => x"8d2d7082",
  1389 => x"2cfc0680",
  1390 => x"da981172",
  1391 => x"109e0671",
  1392 => x"0870722a",
  1393 => x"70830682",
  1394 => x"742b7009",
  1395 => x"7406760c",
  1396 => x"54515657",
  1397 => x"535153a8",
  1398 => x"872d7180",
  1399 => x"dcbc0c02",
  1400 => x"90050d04",
  1401 => x"02fc050d",
  1402 => x"72518071",
  1403 => x"0c800b84",
  1404 => x"120c0284",
  1405 => x"050d0402",
  1406 => x"f0050d75",
  1407 => x"70088412",
  1408 => x"08535353",
  1409 => x"ff547171",
  1410 => x"2ea838a8",
  1411 => x"8d2d8413",
  1412 => x"08708429",
  1413 => x"14881170",
  1414 => x"087081ff",
  1415 => x"06841808",
  1416 => x"81118706",
  1417 => x"841a0c53",
  1418 => x"51555151",
  1419 => x"51a8872d",
  1420 => x"71547380",
  1421 => x"dcbc0c02",
  1422 => x"90050d04",
  1423 => x"02f8050d",
  1424 => x"a88d2de0",
  1425 => x"08708b2a",
  1426 => x"70810651",
  1427 => x"52527080",
  1428 => x"2ea13880",
  1429 => x"ddec0870",
  1430 => x"842980dd",
  1431 => x"f4057381",
  1432 => x"ff06710c",
  1433 => x"515180dd",
  1434 => x"ec088111",
  1435 => x"870680dd",
  1436 => x"ec0c5180",
  1437 => x"0b80de94",
  1438 => x"0ca7ff2d",
  1439 => x"a8872d02",
  1440 => x"88050d04",
  1441 => x"02fc050d",
  1442 => x"a88d2d81",
  1443 => x"0b80de94",
  1444 => x"0ca8872d",
  1445 => x"80de9408",
  1446 => x"5170f938",
  1447 => x"0284050d",
  1448 => x"0402fc05",
  1449 => x"0d80ddec",
  1450 => x"51abe42d",
  1451 => x"ab8b2dac",
  1452 => x"bc51a7fb",
  1453 => x"2d028405",
  1454 => x"0d0480de",
  1455 => x"a00880dc",
  1456 => x"bc0c0402",
  1457 => x"fc050d81",
  1458 => x"0b80dafc",
  1459 => x"0c815185",
  1460 => x"8d2d0284",
  1461 => x"050d0402",
  1462 => x"fc050dad",
  1463 => x"e104a8d8",
  1464 => x"2d80f651",
  1465 => x"aba92d80",
  1466 => x"dcbc08f2",
  1467 => x"3880da51",
  1468 => x"aba92d80",
  1469 => x"dcbc08e6",
  1470 => x"3880dcbc",
  1471 => x"0880dafc",
  1472 => x"0c80dcbc",
  1473 => x"0851858d",
  1474 => x"2d028405",
  1475 => x"0d0402ec",
  1476 => x"050d7654",
  1477 => x"8052870b",
  1478 => x"881580f5",
  1479 => x"2d565374",
  1480 => x"72248338",
  1481 => x"a0537251",
  1482 => x"83842d81",
  1483 => x"128b1580",
  1484 => x"f52d5452",
  1485 => x"727225de",
  1486 => x"38029405",
  1487 => x"0d0402f0",
  1488 => x"050d80de",
  1489 => x"a0085481",
  1490 => x"f92d800b",
  1491 => x"80dea40c",
  1492 => x"7308802e",
  1493 => x"81893882",
  1494 => x"0b80dcd0",
  1495 => x"0c80dea4",
  1496 => x"088f0680",
  1497 => x"dccc0c73",
  1498 => x"08527183",
  1499 => x"2e963871",
  1500 => x"83268938",
  1501 => x"71812eb0",
  1502 => x"38afc804",
  1503 => x"71852ea0",
  1504 => x"38afc804",
  1505 => x"881480f5",
  1506 => x"2d841508",
  1507 => x"80d6f053",
  1508 => x"545286a0",
  1509 => x"2d718429",
  1510 => x"13700852",
  1511 => x"52afcc04",
  1512 => x"7351ae8e",
  1513 => x"2dafc804",
  1514 => x"80daf808",
  1515 => x"8815082c",
  1516 => x"70810651",
  1517 => x"5271802e",
  1518 => x"883880d6",
  1519 => x"f451afc5",
  1520 => x"0480d6f8",
  1521 => x"5186a02d",
  1522 => x"84140851",
  1523 => x"86a02d80",
  1524 => x"dea40881",
  1525 => x"0580dea4",
  1526 => x"0c8c1454",
  1527 => x"aed00402",
  1528 => x"90050d04",
  1529 => x"7180dea0",
  1530 => x"0caebe2d",
  1531 => x"80dea408",
  1532 => x"ff0580de",
  1533 => x"a80c0402",
  1534 => x"e8050d80",
  1535 => x"dea00880",
  1536 => x"deac0857",
  1537 => x"5580f651",
  1538 => x"aba92d80",
  1539 => x"dcbc0881",
  1540 => x"2a708106",
  1541 => x"51527180",
  1542 => x"2ea438b0",
  1543 => x"a104a8d8",
  1544 => x"2d80f651",
  1545 => x"aba92d80",
  1546 => x"dcbc08f2",
  1547 => x"3880dafc",
  1548 => x"08813270",
  1549 => x"80dafc0c",
  1550 => x"70525285",
  1551 => x"8d2d800b",
  1552 => x"80de980c",
  1553 => x"800b80de",
  1554 => x"9c0c80da",
  1555 => x"fc08838d",
  1556 => x"3880da51",
  1557 => x"aba92d80",
  1558 => x"dcbc0880",
  1559 => x"2e8c3880",
  1560 => x"de980881",
  1561 => x"800780de",
  1562 => x"980c80d9",
  1563 => x"51aba92d",
  1564 => x"80dcbc08",
  1565 => x"802e8c38",
  1566 => x"80de9808",
  1567 => x"80c00780",
  1568 => x"de980c81",
  1569 => x"9451aba9",
  1570 => x"2d80dcbc",
  1571 => x"08802e8b",
  1572 => x"3880de98",
  1573 => x"08900780",
  1574 => x"de980c81",
  1575 => x"9151aba9",
  1576 => x"2d80dcbc",
  1577 => x"08802e8b",
  1578 => x"3880de98",
  1579 => x"08a00780",
  1580 => x"de980c81",
  1581 => x"f551aba9",
  1582 => x"2d80dcbc",
  1583 => x"08802e8b",
  1584 => x"3880de98",
  1585 => x"08810780",
  1586 => x"de980c81",
  1587 => x"f251aba9",
  1588 => x"2d80dcbc",
  1589 => x"08802e8b",
  1590 => x"3880de98",
  1591 => x"08820780",
  1592 => x"de980c81",
  1593 => x"eb51aba9",
  1594 => x"2d80dcbc",
  1595 => x"08802e8b",
  1596 => x"3880de98",
  1597 => x"08840780",
  1598 => x"de980c81",
  1599 => x"f451aba9",
  1600 => x"2d80dcbc",
  1601 => x"08802e8b",
  1602 => x"3880de98",
  1603 => x"08880780",
  1604 => x"de980c80",
  1605 => x"d851aba9",
  1606 => x"2d80dcbc",
  1607 => x"08802e8c",
  1608 => x"3880de9c",
  1609 => x"08818007",
  1610 => x"80de9c0c",
  1611 => x"9251aba9",
  1612 => x"2d80dcbc",
  1613 => x"08802e8c",
  1614 => x"3880de9c",
  1615 => x"0880c007",
  1616 => x"80de9c0c",
  1617 => x"9451aba9",
  1618 => x"2d80dcbc",
  1619 => x"08802e8b",
  1620 => x"3880de9c",
  1621 => x"08900780",
  1622 => x"de9c0c91",
  1623 => x"51aba92d",
  1624 => x"80dcbc08",
  1625 => x"802e8b38",
  1626 => x"80de9c08",
  1627 => x"a00780de",
  1628 => x"9c0c9d51",
  1629 => x"aba92d80",
  1630 => x"dcbc0880",
  1631 => x"2e8b3880",
  1632 => x"de9c0881",
  1633 => x"0780de9c",
  1634 => x"0c9b51ab",
  1635 => x"a92d80dc",
  1636 => x"bc08802e",
  1637 => x"8b3880de",
  1638 => x"9c088207",
  1639 => x"80de9c0c",
  1640 => x"9c51aba9",
  1641 => x"2d80dcbc",
  1642 => x"08802e8b",
  1643 => x"3880de9c",
  1644 => x"08840780",
  1645 => x"de9c0ca3",
  1646 => x"51aba92d",
  1647 => x"80dcbc08",
  1648 => x"802e8b38",
  1649 => x"80de9c08",
  1650 => x"880780de",
  1651 => x"9c0c81fd",
  1652 => x"51aba92d",
  1653 => x"81fa51ab",
  1654 => x"a92db9b2",
  1655 => x"0481f551",
  1656 => x"aba92d80",
  1657 => x"dcbc0881",
  1658 => x"2a708106",
  1659 => x"51527180",
  1660 => x"2eb33880",
  1661 => x"dea80852",
  1662 => x"71802e8a",
  1663 => x"38ff1280",
  1664 => x"dea80cb4",
  1665 => x"a50480de",
  1666 => x"a4081080",
  1667 => x"dea40805",
  1668 => x"70842916",
  1669 => x"51528812",
  1670 => x"08802e89",
  1671 => x"38ff5188",
  1672 => x"12085271",
  1673 => x"2d81f251",
  1674 => x"aba92d80",
  1675 => x"dcbc0881",
  1676 => x"2a708106",
  1677 => x"51527180",
  1678 => x"2eb43880",
  1679 => x"dea408ff",
  1680 => x"1180dea8",
  1681 => x"08565353",
  1682 => x"7372258a",
  1683 => x"38811480",
  1684 => x"dea80cb4",
  1685 => x"ee047210",
  1686 => x"13708429",
  1687 => x"16515288",
  1688 => x"1208802e",
  1689 => x"8938fe51",
  1690 => x"88120852",
  1691 => x"712d81fd",
  1692 => x"51aba92d",
  1693 => x"80dcbc08",
  1694 => x"812a7081",
  1695 => x"06515271",
  1696 => x"802eb138",
  1697 => x"80dea808",
  1698 => x"802e8a38",
  1699 => x"800b80de",
  1700 => x"a80cb5b4",
  1701 => x"0480dea4",
  1702 => x"081080de",
  1703 => x"a4080570",
  1704 => x"84291651",
  1705 => x"52881208",
  1706 => x"802e8938",
  1707 => x"fd518812",
  1708 => x"0852712d",
  1709 => x"81fa51ab",
  1710 => x"a92d80dc",
  1711 => x"bc08812a",
  1712 => x"70810651",
  1713 => x"5271802e",
  1714 => x"b13880de",
  1715 => x"a408ff11",
  1716 => x"545280de",
  1717 => x"a8087325",
  1718 => x"89387280",
  1719 => x"dea80cb5",
  1720 => x"fa047110",
  1721 => x"12708429",
  1722 => x"16515288",
  1723 => x"1208802e",
  1724 => x"8938fc51",
  1725 => x"88120852",
  1726 => x"712d80de",
  1727 => x"a8087053",
  1728 => x"5473802e",
  1729 => x"8a388c15",
  1730 => x"ff155555",
  1731 => x"b6810482",
  1732 => x"0b80dcd0",
  1733 => x"0c718f06",
  1734 => x"80dccc0c",
  1735 => x"81eb51ab",
  1736 => x"a92d80dc",
  1737 => x"bc08812a",
  1738 => x"70810651",
  1739 => x"5271802e",
  1740 => x"ad387408",
  1741 => x"852e0981",
  1742 => x"06a43888",
  1743 => x"1580f52d",
  1744 => x"ff055271",
  1745 => x"881681b7",
  1746 => x"2d71982b",
  1747 => x"52718025",
  1748 => x"8838800b",
  1749 => x"881681b7",
  1750 => x"2d7451ae",
  1751 => x"8e2d81f4",
  1752 => x"51aba92d",
  1753 => x"80dcbc08",
  1754 => x"812a7081",
  1755 => x"06515271",
  1756 => x"802eb338",
  1757 => x"7408852e",
  1758 => x"098106aa",
  1759 => x"38881580",
  1760 => x"f52d8105",
  1761 => x"52718816",
  1762 => x"81b72d71",
  1763 => x"81ff068b",
  1764 => x"1680f52d",
  1765 => x"54527272",
  1766 => x"27873872",
  1767 => x"881681b7",
  1768 => x"2d7451ae",
  1769 => x"8e2d80da",
  1770 => x"51aba92d",
  1771 => x"80dcbc08",
  1772 => x"812a7081",
  1773 => x"06515271",
  1774 => x"802e81ad",
  1775 => x"3880dea0",
  1776 => x"0880dea8",
  1777 => x"08555373",
  1778 => x"802e8a38",
  1779 => x"8c13ff15",
  1780 => x"5553b7c7",
  1781 => x"04720852",
  1782 => x"71822ea6",
  1783 => x"38718226",
  1784 => x"89387181",
  1785 => x"2eaa38b8",
  1786 => x"e9047183",
  1787 => x"2eb43871",
  1788 => x"842e0981",
  1789 => x"0680f238",
  1790 => x"88130851",
  1791 => x"afe42db8",
  1792 => x"e90480de",
  1793 => x"a8085188",
  1794 => x"13085271",
  1795 => x"2db8e904",
  1796 => x"810b8814",
  1797 => x"082b80da",
  1798 => x"f8083280",
  1799 => x"daf80cb8",
  1800 => x"bd048813",
  1801 => x"80f52d81",
  1802 => x"058b1480",
  1803 => x"f52d5354",
  1804 => x"71742483",
  1805 => x"38805473",
  1806 => x"881481b7",
  1807 => x"2daebe2d",
  1808 => x"b8e90475",
  1809 => x"08802ea4",
  1810 => x"38750851",
  1811 => x"aba92d80",
  1812 => x"dcbc0881",
  1813 => x"06527180",
  1814 => x"2e8c3880",
  1815 => x"dea80851",
  1816 => x"84160852",
  1817 => x"712d8816",
  1818 => x"5675d838",
  1819 => x"8054800b",
  1820 => x"80dcd00c",
  1821 => x"738f0680",
  1822 => x"dccc0ca0",
  1823 => x"527380de",
  1824 => x"a8082e09",
  1825 => x"81069938",
  1826 => x"80dea408",
  1827 => x"ff057432",
  1828 => x"70098105",
  1829 => x"7072079f",
  1830 => x"2a917131",
  1831 => x"51515353",
  1832 => x"71518384",
  1833 => x"2d811454",
  1834 => x"8e7425c2",
  1835 => x"3880dafc",
  1836 => x"08527180",
  1837 => x"dcbc0c02",
  1838 => x"98050d04",
  1839 => x"02f4050d",
  1840 => x"d45281ff",
  1841 => x"720c7108",
  1842 => x"5381ff72",
  1843 => x"0c72882b",
  1844 => x"83fe8006",
  1845 => x"72087081",
  1846 => x"ff065152",
  1847 => x"5381ff72",
  1848 => x"0c727107",
  1849 => x"882b7208",
  1850 => x"7081ff06",
  1851 => x"51525381",
  1852 => x"ff720c72",
  1853 => x"7107882b",
  1854 => x"72087081",
  1855 => x"ff067207",
  1856 => x"80dcbc0c",
  1857 => x"5253028c",
  1858 => x"050d0402",
  1859 => x"f4050d74",
  1860 => x"767181ff",
  1861 => x"06d40c53",
  1862 => x"5380deb0",
  1863 => x"08853871",
  1864 => x"892b5271",
  1865 => x"982ad40c",
  1866 => x"71902a70",
  1867 => x"81ff06d4",
  1868 => x"0c517188",
  1869 => x"2a7081ff",
  1870 => x"06d40c51",
  1871 => x"7181ff06",
  1872 => x"d40c7290",
  1873 => x"2a7081ff",
  1874 => x"06d40c51",
  1875 => x"d4087081",
  1876 => x"ff065151",
  1877 => x"82b8bf52",
  1878 => x"7081ff2e",
  1879 => x"09810694",
  1880 => x"3881ff0b",
  1881 => x"d40cd408",
  1882 => x"7081ff06",
  1883 => x"ff145451",
  1884 => x"5171e538",
  1885 => x"7080dcbc",
  1886 => x"0c028c05",
  1887 => x"0d0402fc",
  1888 => x"050d81c7",
  1889 => x"5181ff0b",
  1890 => x"d40cff11",
  1891 => x"51708025",
  1892 => x"f4380284",
  1893 => x"050d0402",
  1894 => x"f4050d81",
  1895 => x"ff0bd40c",
  1896 => x"93538052",
  1897 => x"87fc80c1",
  1898 => x"51ba8b2d",
  1899 => x"80dcbc08",
  1900 => x"8b3881ff",
  1901 => x"0bd40c81",
  1902 => x"53bbc504",
  1903 => x"bafe2dff",
  1904 => x"135372de",
  1905 => x"387280dc",
  1906 => x"bc0c028c",
  1907 => x"050d0402",
  1908 => x"ec050d81",
  1909 => x"0b80deb0",
  1910 => x"0c8454d0",
  1911 => x"08708f2a",
  1912 => x"70810651",
  1913 => x"515372f3",
  1914 => x"3872d00c",
  1915 => x"bafe2d80",
  1916 => x"d6fc5186",
  1917 => x"a02dd008",
  1918 => x"708f2a70",
  1919 => x"81065151",
  1920 => x"5372f338",
  1921 => x"810bd00c",
  1922 => x"b1538052",
  1923 => x"84d480c0",
  1924 => x"51ba8b2d",
  1925 => x"80dcbc08",
  1926 => x"812e9338",
  1927 => x"72822ebf",
  1928 => x"38ff1353",
  1929 => x"72e438ff",
  1930 => x"145473ff",
  1931 => x"ae38bafe",
  1932 => x"2d83aa52",
  1933 => x"849c80c8",
  1934 => x"51ba8b2d",
  1935 => x"80dcbc08",
  1936 => x"812e0981",
  1937 => x"069338b9",
  1938 => x"bc2d80dc",
  1939 => x"bc0883ff",
  1940 => x"ff065372",
  1941 => x"83aa2e9f",
  1942 => x"38bb972d",
  1943 => x"bcf20480",
  1944 => x"d7885186",
  1945 => x"a02d8053",
  1946 => x"bec70480",
  1947 => x"d7a05186",
  1948 => x"a02d8054",
  1949 => x"be980481",
  1950 => x"ff0bd40c",
  1951 => x"b154bafe",
  1952 => x"2d8fcf53",
  1953 => x"805287fc",
  1954 => x"80f751ba",
  1955 => x"8b2d80dc",
  1956 => x"bc085580",
  1957 => x"dcbc0881",
  1958 => x"2e098106",
  1959 => x"9c3881ff",
  1960 => x"0bd40c82",
  1961 => x"0a52849c",
  1962 => x"80e951ba",
  1963 => x"8b2d80dc",
  1964 => x"bc08802e",
  1965 => x"8d38bafe",
  1966 => x"2dff1353",
  1967 => x"72c638be",
  1968 => x"8b0481ff",
  1969 => x"0bd40c80",
  1970 => x"dcbc0852",
  1971 => x"87fc80fa",
  1972 => x"51ba8b2d",
  1973 => x"80dcbc08",
  1974 => x"b23881ff",
  1975 => x"0bd40cd4",
  1976 => x"085381ff",
  1977 => x"0bd40c81",
  1978 => x"ff0bd40c",
  1979 => x"81ff0bd4",
  1980 => x"0c81ff0b",
  1981 => x"d40c7286",
  1982 => x"2a708106",
  1983 => x"76565153",
  1984 => x"72963880",
  1985 => x"dcbc0854",
  1986 => x"be980473",
  1987 => x"822efedb",
  1988 => x"38ff1454",
  1989 => x"73fee738",
  1990 => x"7380deb0",
  1991 => x"0c738b38",
  1992 => x"815287fc",
  1993 => x"80d051ba",
  1994 => x"8b2d81ff",
  1995 => x"0bd40cd0",
  1996 => x"08708f2a",
  1997 => x"70810651",
  1998 => x"515372f3",
  1999 => x"3872d00c",
  2000 => x"81ff0bd4",
  2001 => x"0c815372",
  2002 => x"80dcbc0c",
  2003 => x"0294050d",
  2004 => x"0402e805",
  2005 => x"0d785580",
  2006 => x"5681ff0b",
  2007 => x"d40cd008",
  2008 => x"708f2a70",
  2009 => x"81065151",
  2010 => x"5372f338",
  2011 => x"82810bd0",
  2012 => x"0c81ff0b",
  2013 => x"d40c7752",
  2014 => x"87fc80d1",
  2015 => x"51ba8b2d",
  2016 => x"80dbc6df",
  2017 => x"5480dcbc",
  2018 => x"08802e8b",
  2019 => x"3880d7c0",
  2020 => x"5186a02d",
  2021 => x"bfeb0481",
  2022 => x"ff0bd40c",
  2023 => x"d4087081",
  2024 => x"ff065153",
  2025 => x"7281fe2e",
  2026 => x"0981069e",
  2027 => x"3880ff53",
  2028 => x"b9bc2d80",
  2029 => x"dcbc0875",
  2030 => x"70840557",
  2031 => x"0cff1353",
  2032 => x"728025ec",
  2033 => x"388156bf",
  2034 => x"d004ff14",
  2035 => x"5473c838",
  2036 => x"81ff0bd4",
  2037 => x"0c81ff0b",
  2038 => x"d40cd008",
  2039 => x"708f2a70",
  2040 => x"81065151",
  2041 => x"5372f338",
  2042 => x"72d00c75",
  2043 => x"80dcbc0c",
  2044 => x"0298050d",
  2045 => x"0402e805",
  2046 => x"0d77797b",
  2047 => x"58555580",
  2048 => x"53727625",
  2049 => x"a5387470",
  2050 => x"81055680",
  2051 => x"f52d7470",
  2052 => x"81055680",
  2053 => x"f52d5252",
  2054 => x"71712e87",
  2055 => x"38815180",
  2056 => x"c0ac0481",
  2057 => x"135380c0",
  2058 => x"81048051",
  2059 => x"7080dcbc",
  2060 => x"0c029805",
  2061 => x"0d0402ec",
  2062 => x"050d7655",
  2063 => x"74802e80",
  2064 => x"c4389a15",
  2065 => x"80e02d51",
  2066 => x"80cee42d",
  2067 => x"80dcbc08",
  2068 => x"80dcbc08",
  2069 => x"80e4e40c",
  2070 => x"80dcbc08",
  2071 => x"545480e4",
  2072 => x"c008802e",
  2073 => x"9b389415",
  2074 => x"80e02d51",
  2075 => x"80cee42d",
  2076 => x"80dcbc08",
  2077 => x"902b83ff",
  2078 => x"f00a0670",
  2079 => x"75075153",
  2080 => x"7280e4e4",
  2081 => x"0c80e4e4",
  2082 => x"08537280",
  2083 => x"2e9e3880",
  2084 => x"e4b808fe",
  2085 => x"14712980",
  2086 => x"e4cc0805",
  2087 => x"80e4e80c",
  2088 => x"70842b80",
  2089 => x"e4c40c54",
  2090 => x"80c1db04",
  2091 => x"80e4d008",
  2092 => x"80e4e40c",
  2093 => x"80e4d408",
  2094 => x"80e4e80c",
  2095 => x"80e4c008",
  2096 => x"802e8c38",
  2097 => x"80e4b808",
  2098 => x"842b5380",
  2099 => x"c1d60480",
  2100 => x"e4d80884",
  2101 => x"2b537280",
  2102 => x"e4c40c02",
  2103 => x"94050d04",
  2104 => x"02d8050d",
  2105 => x"800b80e4",
  2106 => x"c00c8454",
  2107 => x"bbcf2d80",
  2108 => x"dcbc0880",
  2109 => x"2e983880",
  2110 => x"deb45280",
  2111 => x"51bed12d",
  2112 => x"80dcbc08",
  2113 => x"802e8738",
  2114 => x"fe5480c2",
  2115 => x"9604ff14",
  2116 => x"54738024",
  2117 => x"d738738e",
  2118 => x"3880d7d0",
  2119 => x"5186a02d",
  2120 => x"735580c7",
  2121 => x"f4048056",
  2122 => x"810b80e4",
  2123 => x"ec0c8853",
  2124 => x"80d7e452",
  2125 => x"80deea51",
  2126 => x"bff52d80",
  2127 => x"dcbc0876",
  2128 => x"2e098106",
  2129 => x"893880dc",
  2130 => x"bc0880e4",
  2131 => x"ec0c8853",
  2132 => x"80d7f052",
  2133 => x"80df8651",
  2134 => x"bff52d80",
  2135 => x"dcbc0889",
  2136 => x"3880dcbc",
  2137 => x"0880e4ec",
  2138 => x"0c80e4ec",
  2139 => x"08802e81",
  2140 => x"843880e1",
  2141 => x"fa0b80f5",
  2142 => x"2d80e1fb",
  2143 => x"0b80f52d",
  2144 => x"71982b71",
  2145 => x"902b0780",
  2146 => x"e1fc0b80",
  2147 => x"f52d7088",
  2148 => x"2b720780",
  2149 => x"e1fd0b80",
  2150 => x"f52d7107",
  2151 => x"80e2b20b",
  2152 => x"80f52d80",
  2153 => x"e2b30b80",
  2154 => x"f52d7188",
  2155 => x"2b07535f",
  2156 => x"54525a56",
  2157 => x"57557381",
  2158 => x"abaa2e09",
  2159 => x"81069038",
  2160 => x"755180ce",
  2161 => x"b32d80dc",
  2162 => x"bc085680",
  2163 => x"c3de0473",
  2164 => x"82d4d52e",
  2165 => x"893880d7",
  2166 => x"fc5180c4",
  2167 => x"ab0480de",
  2168 => x"b4527551",
  2169 => x"bed12d80",
  2170 => x"dcbc0855",
  2171 => x"80dcbc08",
  2172 => x"802e8480",
  2173 => x"38885380",
  2174 => x"d7f05280",
  2175 => x"df8651bf",
  2176 => x"f52d80dc",
  2177 => x"bc088b38",
  2178 => x"810b80e4",
  2179 => x"c00c80c4",
  2180 => x"b2048853",
  2181 => x"80d7e452",
  2182 => x"80deea51",
  2183 => x"bff52d80",
  2184 => x"dcbc0880",
  2185 => x"2e8c3880",
  2186 => x"d8905186",
  2187 => x"a02d80c5",
  2188 => x"910480e2",
  2189 => x"b20b80f5",
  2190 => x"2d547380",
  2191 => x"d52e0981",
  2192 => x"0680ce38",
  2193 => x"80e2b30b",
  2194 => x"80f52d54",
  2195 => x"7381aa2e",
  2196 => x"098106bd",
  2197 => x"38800b80",
  2198 => x"deb40b80",
  2199 => x"f52d5654",
  2200 => x"7481e92e",
  2201 => x"83388154",
  2202 => x"7481eb2e",
  2203 => x"8c388055",
  2204 => x"73752e09",
  2205 => x"810682fc",
  2206 => x"3880debf",
  2207 => x"0b80f52d",
  2208 => x"55748e38",
  2209 => x"80dec00b",
  2210 => x"80f52d54",
  2211 => x"73822e87",
  2212 => x"38805580",
  2213 => x"c7f40480",
  2214 => x"dec10b80",
  2215 => x"f52d7080",
  2216 => x"e4b80cff",
  2217 => x"0580e4bc",
  2218 => x"0c80dec2",
  2219 => x"0b80f52d",
  2220 => x"80dec30b",
  2221 => x"80f52d58",
  2222 => x"76057782",
  2223 => x"80290570",
  2224 => x"80e4c80c",
  2225 => x"80dec40b",
  2226 => x"80f52d70",
  2227 => x"80e4dc0c",
  2228 => x"80e4c008",
  2229 => x"59575876",
  2230 => x"802e81b8",
  2231 => x"38885380",
  2232 => x"d7f05280",
  2233 => x"df8651bf",
  2234 => x"f52d80dc",
  2235 => x"bc088284",
  2236 => x"3880e4b8",
  2237 => x"0870842b",
  2238 => x"80e4c40c",
  2239 => x"7080e4d8",
  2240 => x"0c80ded9",
  2241 => x"0b80f52d",
  2242 => x"80ded80b",
  2243 => x"80f52d71",
  2244 => x"82802905",
  2245 => x"80deda0b",
  2246 => x"80f52d70",
  2247 => x"84808029",
  2248 => x"1280dedb",
  2249 => x"0b80f52d",
  2250 => x"7081800a",
  2251 => x"29127080",
  2252 => x"e4e00c80",
  2253 => x"e4dc0871",
  2254 => x"2980e4c8",
  2255 => x"08057080",
  2256 => x"e4cc0c80",
  2257 => x"dee10b80",
  2258 => x"f52d80de",
  2259 => x"e00b80f5",
  2260 => x"2d718280",
  2261 => x"290580de",
  2262 => x"e20b80f5",
  2263 => x"2d708480",
  2264 => x"80291280",
  2265 => x"dee30b80",
  2266 => x"f52d7098",
  2267 => x"2b81f00a",
  2268 => x"06720570",
  2269 => x"80e4d00c",
  2270 => x"fe117e29",
  2271 => x"770580e4",
  2272 => x"d40c5259",
  2273 => x"5243545e",
  2274 => x"51525952",
  2275 => x"5d575957",
  2276 => x"80c7ec04",
  2277 => x"80dec60b",
  2278 => x"80f52d80",
  2279 => x"dec50b80",
  2280 => x"f52d7182",
  2281 => x"80290570",
  2282 => x"80e4c40c",
  2283 => x"70a02983",
  2284 => x"ff057089",
  2285 => x"2a7080e4",
  2286 => x"d80c80de",
  2287 => x"cb0b80f5",
  2288 => x"2d80deca",
  2289 => x"0b80f52d",
  2290 => x"71828029",
  2291 => x"057080e4",
  2292 => x"e00c7b71",
  2293 => x"291e7080",
  2294 => x"e4d40c7d",
  2295 => x"80e4d00c",
  2296 => x"730580e4",
  2297 => x"cc0c555e",
  2298 => x"51515555",
  2299 => x"805180c0",
  2300 => x"b62d8155",
  2301 => x"7480dcbc",
  2302 => x"0c02a805",
  2303 => x"0d0402ec",
  2304 => x"050d7670",
  2305 => x"872c7180",
  2306 => x"ff065556",
  2307 => x"5480e4c0",
  2308 => x"088a3873",
  2309 => x"882c7481",
  2310 => x"ff065455",
  2311 => x"80deb452",
  2312 => x"80e4c808",
  2313 => x"1551bed1",
  2314 => x"2d80dcbc",
  2315 => x"085480dc",
  2316 => x"bc08802e",
  2317 => x"bb3880e4",
  2318 => x"c008802e",
  2319 => x"9c387284",
  2320 => x"2980deb4",
  2321 => x"05700852",
  2322 => x"5380ceb3",
  2323 => x"2d80dcbc",
  2324 => x"08f00a06",
  2325 => x"5380c8ee",
  2326 => x"04721080",
  2327 => x"deb40570",
  2328 => x"80e02d52",
  2329 => x"5380cee4",
  2330 => x"2d80dcbc",
  2331 => x"08537254",
  2332 => x"7380dcbc",
  2333 => x"0c029405",
  2334 => x"0d0402e0",
  2335 => x"050d7970",
  2336 => x"842c80e4",
  2337 => x"e8080571",
  2338 => x"8f065255",
  2339 => x"53728a38",
  2340 => x"80deb452",
  2341 => x"7351bed1",
  2342 => x"2d72a029",
  2343 => x"80deb405",
  2344 => x"54807480",
  2345 => x"f52d5653",
  2346 => x"74732e83",
  2347 => x"38815374",
  2348 => x"81e52e81",
  2349 => x"f5388170",
  2350 => x"74065458",
  2351 => x"72802e81",
  2352 => x"e9388b14",
  2353 => x"80f52d70",
  2354 => x"832a7906",
  2355 => x"5856769c",
  2356 => x"3880db80",
  2357 => x"08537289",
  2358 => x"387280e2",
  2359 => x"b40b81b7",
  2360 => x"2d7680db",
  2361 => x"800c7353",
  2362 => x"80cbac04",
  2363 => x"758f2e09",
  2364 => x"810681b6",
  2365 => x"38749f06",
  2366 => x"8d2980e2",
  2367 => x"a7115153",
  2368 => x"811480f5",
  2369 => x"2d737081",
  2370 => x"055581b7",
  2371 => x"2d831480",
  2372 => x"f52d7370",
  2373 => x"81055581",
  2374 => x"b72d8514",
  2375 => x"80f52d73",
  2376 => x"70810555",
  2377 => x"81b72d87",
  2378 => x"1480f52d",
  2379 => x"73708105",
  2380 => x"5581b72d",
  2381 => x"891480f5",
  2382 => x"2d737081",
  2383 => x"055581b7",
  2384 => x"2d8e1480",
  2385 => x"f52d7370",
  2386 => x"81055581",
  2387 => x"b72d9014",
  2388 => x"80f52d73",
  2389 => x"70810555",
  2390 => x"81b72d92",
  2391 => x"1480f52d",
  2392 => x"73708105",
  2393 => x"5581b72d",
  2394 => x"941480f5",
  2395 => x"2d737081",
  2396 => x"055581b7",
  2397 => x"2d961480",
  2398 => x"f52d7370",
  2399 => x"81055581",
  2400 => x"b72d9814",
  2401 => x"80f52d73",
  2402 => x"70810555",
  2403 => x"81b72d9c",
  2404 => x"1480f52d",
  2405 => x"73708105",
  2406 => x"5581b72d",
  2407 => x"9e1480f5",
  2408 => x"2d7381b7",
  2409 => x"2d7780db",
  2410 => x"800c8053",
  2411 => x"7280dcbc",
  2412 => x"0c02a005",
  2413 => x"0d0402cc",
  2414 => x"050d7e60",
  2415 => x"5e5a800b",
  2416 => x"80e4e408",
  2417 => x"80e4e808",
  2418 => x"595c5680",
  2419 => x"5880e4c4",
  2420 => x"08782e81",
  2421 => x"bc38778f",
  2422 => x"06a01757",
  2423 => x"54739138",
  2424 => x"80deb452",
  2425 => x"76518117",
  2426 => x"57bed12d",
  2427 => x"80deb456",
  2428 => x"807680f5",
  2429 => x"2d565474",
  2430 => x"742e8338",
  2431 => x"81547481",
  2432 => x"e52e8181",
  2433 => x"38817075",
  2434 => x"06555c73",
  2435 => x"802e80f5",
  2436 => x"388b1680",
  2437 => x"f52d9806",
  2438 => x"597880e9",
  2439 => x"388b537c",
  2440 => x"527551bf",
  2441 => x"f52d80dc",
  2442 => x"bc0880d9",
  2443 => x"389c1608",
  2444 => x"5180ceb3",
  2445 => x"2d80dcbc",
  2446 => x"08841b0c",
  2447 => x"9a1680e0",
  2448 => x"2d5180ce",
  2449 => x"e42d80dc",
  2450 => x"bc0880dc",
  2451 => x"bc08881c",
  2452 => x"0c80dcbc",
  2453 => x"08555580",
  2454 => x"e4c00880",
  2455 => x"2e9a3894",
  2456 => x"1680e02d",
  2457 => x"5180cee4",
  2458 => x"2d80dcbc",
  2459 => x"08902b83",
  2460 => x"fff00a06",
  2461 => x"70165154",
  2462 => x"73881b0c",
  2463 => x"787a0c7b",
  2464 => x"5480cdcf",
  2465 => x"04811858",
  2466 => x"80e4c408",
  2467 => x"7826fec6",
  2468 => x"3880e4c0",
  2469 => x"08802eb5",
  2470 => x"387a5180",
  2471 => x"c7fe2d80",
  2472 => x"dcbc0880",
  2473 => x"dcbc0880",
  2474 => x"fffffff8",
  2475 => x"06555b73",
  2476 => x"80ffffff",
  2477 => x"f82e9638",
  2478 => x"80dcbc08",
  2479 => x"fe0580e4",
  2480 => x"b8082980",
  2481 => x"e4cc0805",
  2482 => x"5780cbcb",
  2483 => x"04805473",
  2484 => x"80dcbc0c",
  2485 => x"02b4050d",
  2486 => x"0402f405",
  2487 => x"0d747008",
  2488 => x"8105710c",
  2489 => x"700880e4",
  2490 => x"bc080653",
  2491 => x"53719038",
  2492 => x"88130851",
  2493 => x"80c7fe2d",
  2494 => x"80dcbc08",
  2495 => x"88140c81",
  2496 => x"0b80dcbc",
  2497 => x"0c028c05",
  2498 => x"0d0402f0",
  2499 => x"050d7588",
  2500 => x"1108fe05",
  2501 => x"80e4b808",
  2502 => x"2980e4cc",
  2503 => x"08117208",
  2504 => x"80e4bc08",
  2505 => x"06057955",
  2506 => x"535454be",
  2507 => x"d12d0290",
  2508 => x"050d0402",
  2509 => x"f4050d74",
  2510 => x"70882a83",
  2511 => x"fe800670",
  2512 => x"72982a07",
  2513 => x"72882b87",
  2514 => x"fc808006",
  2515 => x"73982b81",
  2516 => x"f00a0671",
  2517 => x"73070780",
  2518 => x"dcbc0c56",
  2519 => x"51535102",
  2520 => x"8c050d04",
  2521 => x"02f8050d",
  2522 => x"028e0580",
  2523 => x"f52d7488",
  2524 => x"2b077083",
  2525 => x"ffff0680",
  2526 => x"dcbc0c51",
  2527 => x"0288050d",
  2528 => x"0402f405",
  2529 => x"0d747678",
  2530 => x"53545280",
  2531 => x"71259738",
  2532 => x"72708105",
  2533 => x"5480f52d",
  2534 => x"72708105",
  2535 => x"5481b72d",
  2536 => x"ff115170",
  2537 => x"eb388072",
  2538 => x"81b72d02",
  2539 => x"8c050d04",
  2540 => x"02e8050d",
  2541 => x"77568070",
  2542 => x"56547376",
  2543 => x"24b73880",
  2544 => x"e4c40874",
  2545 => x"2eaf3873",
  2546 => x"5180c8fa",
  2547 => x"2d80dcbc",
  2548 => x"0880dcbc",
  2549 => x"08098105",
  2550 => x"7080dcbc",
  2551 => x"08079f2a",
  2552 => x"77058117",
  2553 => x"57575353",
  2554 => x"74762489",
  2555 => x"3880e4c4",
  2556 => x"087426d3",
  2557 => x"387280dc",
  2558 => x"bc0c0298",
  2559 => x"050d0402",
  2560 => x"f0050d80",
  2561 => x"dcb80816",
  2562 => x"5180cfb0",
  2563 => x"2d80dcbc",
  2564 => x"08802ea0",
  2565 => x"388b5380",
  2566 => x"dcbc0852",
  2567 => x"80e2b451",
  2568 => x"80cf812d",
  2569 => x"80e4f008",
  2570 => x"5473802e",
  2571 => x"873880e2",
  2572 => x"b451732d",
  2573 => x"0290050d",
  2574 => x"0402dc05",
  2575 => x"0d80705a",
  2576 => x"557480dc",
  2577 => x"b80825b5",
  2578 => x"3880e4c4",
  2579 => x"08752ead",
  2580 => x"38785180",
  2581 => x"c8fa2d80",
  2582 => x"dcbc0809",
  2583 => x"81057080",
  2584 => x"dcbc0807",
  2585 => x"9f2a7605",
  2586 => x"811b5b56",
  2587 => x"547480dc",
  2588 => x"b8082589",
  2589 => x"3880e4c4",
  2590 => x"087926d5",
  2591 => x"38805578",
  2592 => x"80e4c408",
  2593 => x"2781e438",
  2594 => x"785180c8",
  2595 => x"fa2d80dc",
  2596 => x"bc08802e",
  2597 => x"81b43880",
  2598 => x"dcbc088b",
  2599 => x"0580f52d",
  2600 => x"70842a70",
  2601 => x"81067710",
  2602 => x"78842b80",
  2603 => x"e2b40b80",
  2604 => x"f52d5c5c",
  2605 => x"53515556",
  2606 => x"73802e80",
  2607 => x"ce387416",
  2608 => x"822b80d3",
  2609 => x"8f0b80db",
  2610 => x"8c120c54",
  2611 => x"77753110",
  2612 => x"80e4f411",
  2613 => x"55569074",
  2614 => x"70810556",
  2615 => x"81b72da0",
  2616 => x"7481b72d",
  2617 => x"7681ff06",
  2618 => x"81165854",
  2619 => x"73802e8b",
  2620 => x"389c5380",
  2621 => x"e2b45280",
  2622 => x"d282048b",
  2623 => x"5380dcbc",
  2624 => x"085280e4",
  2625 => x"f6165180",
  2626 => x"d2c00474",
  2627 => x"16822b80",
  2628 => x"cfff0b80",
  2629 => x"db8c120c",
  2630 => x"547681ff",
  2631 => x"06811658",
  2632 => x"5473802e",
  2633 => x"8b389c53",
  2634 => x"80e2b452",
  2635 => x"80d2b704",
  2636 => x"8b5380dc",
  2637 => x"bc085277",
  2638 => x"75311080",
  2639 => x"e4f40551",
  2640 => x"765580cf",
  2641 => x"812d80d2",
  2642 => x"df047490",
  2643 => x"29753170",
  2644 => x"1080e4f4",
  2645 => x"05515480",
  2646 => x"dcbc0874",
  2647 => x"81b72d81",
  2648 => x"1959748b",
  2649 => x"24a43880",
  2650 => x"d0ff0474",
  2651 => x"90297531",
  2652 => x"701080e4",
  2653 => x"f4058c77",
  2654 => x"31575154",
  2655 => x"807481b7",
  2656 => x"2d9e14ff",
  2657 => x"16565474",
  2658 => x"f33802a4",
  2659 => x"050d0402",
  2660 => x"fc050d80",
  2661 => x"dcb80813",
  2662 => x"5180cfb0",
  2663 => x"2d80dcbc",
  2664 => x"08802e8a",
  2665 => x"3880dcbc",
  2666 => x"085180c0",
  2667 => x"b62d800b",
  2668 => x"80dcb80c",
  2669 => x"80d0b92d",
  2670 => x"aebe2d02",
  2671 => x"84050d04",
  2672 => x"02fc050d",
  2673 => x"725170fd",
  2674 => x"2eb23870",
  2675 => x"fd248b38",
  2676 => x"70fc2e80",
  2677 => x"d03880d4",
  2678 => x"af0470fe",
  2679 => x"2eb93870",
  2680 => x"ff2e0981",
  2681 => x"0680c838",
  2682 => x"80dcb808",
  2683 => x"5170802e",
  2684 => x"be38ff11",
  2685 => x"80dcb80c",
  2686 => x"80d4af04",
  2687 => x"80dcb808",
  2688 => x"f0057080",
  2689 => x"dcb80c51",
  2690 => x"708025a3",
  2691 => x"38800b80",
  2692 => x"dcb80c80",
  2693 => x"d4af0480",
  2694 => x"dcb80881",
  2695 => x"0580dcb8",
  2696 => x"0c80d4af",
  2697 => x"0480dcb8",
  2698 => x"08900580",
  2699 => x"dcb80c80",
  2700 => x"d0b92dae",
  2701 => x"be2d0284",
  2702 => x"050d0402",
  2703 => x"fc050d80",
  2704 => x"0b80dcb8",
  2705 => x"0c80d0b9",
  2706 => x"2dadba2d",
  2707 => x"80dcbc08",
  2708 => x"80dca80c",
  2709 => x"80db8451",
  2710 => x"afe42d02",
  2711 => x"84050d04",
  2712 => x"7180e4f0",
  2713 => x"0c040000",
  2714 => x"00ffffff",
  2715 => x"ff00ffff",
  2716 => x"ffff00ff",
  2717 => x"ffffff00",
  2718 => x"30313233",
  2719 => x"34353637",
  2720 => x"38394142",
  2721 => x"43444546",
  2722 => x"00000000",
  2723 => x"44656275",
  2724 => x"67000000",
  2725 => x"52657365",
  2726 => x"74000000",
  2727 => x"5363616e",
  2728 => x"6c696e65",
  2729 => x"73000000",
  2730 => x"50414c20",
  2731 => x"2f204e54",
  2732 => x"53430000",
  2733 => x"436f6c6f",
  2734 => x"72000000",
  2735 => x"44696666",
  2736 => x"6963756c",
  2737 => x"74792041",
  2738 => x"00000000",
  2739 => x"44696666",
  2740 => x"6963756c",
  2741 => x"74792042",
  2742 => x"00000000",
  2743 => x"2a537570",
  2744 => x"65726368",
  2745 => x"69702069",
  2746 => x"6e206361",
  2747 => x"72747269",
  2748 => x"64676500",
  2749 => x"2a42616e",
  2750 => x"6b204530",
  2751 => x"00000000",
  2752 => x"2a42616e",
  2753 => x"6b204537",
  2754 => x"00000000",
  2755 => x"53656c65",
  2756 => x"63740000",
  2757 => x"53746172",
  2758 => x"74000000",
  2759 => x"4c6f6164",
  2760 => x"20524f4d",
  2761 => x"20100000",
  2762 => x"45786974",
  2763 => x"00000000",
  2764 => x"524f4d20",
  2765 => x"6c6f6164",
  2766 => x"696e6720",
  2767 => x"6661696c",
  2768 => x"65640000",
  2769 => x"4f4b0000",
  2770 => x"496e6974",
  2771 => x"69616c69",
  2772 => x"7a696e67",
  2773 => x"20534420",
  2774 => x"63617264",
  2775 => x"0a000000",
  2776 => x"436f6c6c",
  2777 => x"6563746f",
  2778 => x"72566973",
  2779 => x"696f6e00",
  2780 => x"16200000",
  2781 => x"14200000",
  2782 => x"15200000",
  2783 => x"53442069",
  2784 => x"6e69742e",
  2785 => x"2e2e0a00",
  2786 => x"53442063",
  2787 => x"61726420",
  2788 => x"72657365",
  2789 => x"74206661",
  2790 => x"696c6564",
  2791 => x"210a0000",
  2792 => x"53444843",
  2793 => x"20657272",
  2794 => x"6f72210a",
  2795 => x"00000000",
  2796 => x"57726974",
  2797 => x"65206661",
  2798 => x"696c6564",
  2799 => x"0a000000",
  2800 => x"52656164",
  2801 => x"20666169",
  2802 => x"6c65640a",
  2803 => x"00000000",
  2804 => x"43617264",
  2805 => x"20696e69",
  2806 => x"74206661",
  2807 => x"696c6564",
  2808 => x"0a000000",
  2809 => x"46415431",
  2810 => x"36202020",
  2811 => x"00000000",
  2812 => x"46415433",
  2813 => x"32202020",
  2814 => x"00000000",
  2815 => x"4e6f2070",
  2816 => x"61727469",
  2817 => x"74696f6e",
  2818 => x"20736967",
  2819 => x"0a000000",
  2820 => x"42616420",
  2821 => x"70617274",
  2822 => x"0a000000",
  2823 => x"4261636b",
  2824 => x"00000000",
  2825 => x"00000002",
  2826 => x"00002a78",
  2827 => x"00002ea8",
  2828 => x"00000002",
  2829 => x"00002e64",
  2830 => x"000012e6",
  2831 => x"00000002",
  2832 => x"00002a8c",
  2833 => x"00001276",
  2834 => x"00000002",
  2835 => x"00002a94",
  2836 => x"0000035a",
  2837 => x"00000001",
  2838 => x"00002a9c",
  2839 => x"00000000",
  2840 => x"00000001",
  2841 => x"00002aa8",
  2842 => x"00000001",
  2843 => x"00000001",
  2844 => x"00002ab4",
  2845 => x"00000002",
  2846 => x"00000001",
  2847 => x"00002abc",
  2848 => x"00000003",
  2849 => x"00000001",
  2850 => x"00002acc",
  2851 => x"00000004",
  2852 => x"00000001",
  2853 => x"00002adc",
  2854 => x"00000005",
  2855 => x"00000001",
  2856 => x"00002af4",
  2857 => x"00000008",
  2858 => x"00000001",
  2859 => x"00002b00",
  2860 => x"00000009",
  2861 => x"00000002",
  2862 => x"00002b0c",
  2863 => x"0000036e",
  2864 => x"00000002",
  2865 => x"00002b14",
  2866 => x"00000a3f",
  2867 => x"00000002",
  2868 => x"00002b1c",
  2869 => x"00002a3b",
  2870 => x"00000002",
  2871 => x"00002b28",
  2872 => x"000016d7",
  2873 => x"00000000",
  2874 => x"00000000",
  2875 => x"00000000",
  2876 => x"00000004",
  2877 => x"00002b30",
  2878 => x"00002cf0",
  2879 => x"00000004",
  2880 => x"00002b44",
  2881 => x"00002c30",
  2882 => x"00000000",
  2883 => x"00000000",
  2884 => x"00000000",
  2885 => x"00000000",
  2886 => x"00000000",
  2887 => x"00000000",
  2888 => x"00000000",
  2889 => x"00000000",
  2890 => x"00000000",
  2891 => x"00000000",
  2892 => x"00000000",
  2893 => x"00000000",
  2894 => x"00000000",
  2895 => x"00000000",
  2896 => x"00000000",
  2897 => x"00000000",
  2898 => x"00000000",
  2899 => x"00000000",
  2900 => x"00000000",
  2901 => x"00000000",
  2902 => x"76f55a1c",
  2903 => x"f21c1c1c",
  2904 => x"1c1c1c1c",
  2905 => x"00000000",
  2906 => x"00000fff",
  2907 => x"00000fff",
  2908 => x"00000000",
  2909 => x"00000000",
  2910 => x"00000006",
  2911 => x"00000000",
  2912 => x"00000000",
  2913 => x"00000002",
  2914 => x"00003274",
  2915 => x"000027ff",
  2916 => x"00000002",
  2917 => x"00003292",
  2918 => x"000027ff",
  2919 => x"00000002",
  2920 => x"000032b0",
  2921 => x"000027ff",
  2922 => x"00000002",
  2923 => x"000032ce",
  2924 => x"000027ff",
  2925 => x"00000002",
  2926 => x"000032ec",
  2927 => x"000027ff",
  2928 => x"00000002",
  2929 => x"0000330a",
  2930 => x"000027ff",
  2931 => x"00000002",
  2932 => x"00003328",
  2933 => x"000027ff",
  2934 => x"00000002",
  2935 => x"00003346",
  2936 => x"000027ff",
  2937 => x"00000002",
  2938 => x"00003364",
  2939 => x"000027ff",
  2940 => x"00000002",
  2941 => x"00003382",
  2942 => x"000027ff",
  2943 => x"00000002",
  2944 => x"000033a0",
  2945 => x"000027ff",
  2946 => x"00000002",
  2947 => x"000033be",
  2948 => x"000027ff",
  2949 => x"00000002",
  2950 => x"000033dc",
  2951 => x"000027ff",
  2952 => x"00000004",
  2953 => x"00002c1c",
  2954 => x"00000000",
  2955 => x"00000000",
  2956 => x"00000000",
  2957 => x"000029c0",
  2958 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

