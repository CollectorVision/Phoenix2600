-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80de",
     9 => x"f8080b0b",
    10 => x"80defc08",
    11 => x"0b0b80df",
    12 => x"80080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"df800c0b",
    16 => x"0b80defc",
    17 => x"0c0b0b80",
    18 => x"def80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d6e4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80def870",
    57 => x"80e9b027",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a6d9",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80df",
    65 => x"880c9f0b",
    66 => x"80df8c0c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"df8c08ff",
    70 => x"0580df8c",
    71 => x"0c80df8c",
    72 => x"088025e8",
    73 => x"3880df88",
    74 => x"08ff0580",
    75 => x"df880c80",
    76 => x"df880880",
    77 => x"25d03880",
    78 => x"0b80df8c",
    79 => x"0c800b80",
    80 => x"df880c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80df8808",
   100 => x"25913882",
   101 => x"c82d80df",
   102 => x"8808ff05",
   103 => x"80df880c",
   104 => x"838a0480",
   105 => x"df880880",
   106 => x"df8c0853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80df8808",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"df8c0881",
   116 => x"0580df8c",
   117 => x"0c80df8c",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80df8c",
   121 => x"0c80df88",
   122 => x"08810580",
   123 => x"df880c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480df",
   128 => x"8c088105",
   129 => x"80df8c0c",
   130 => x"80df8c08",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80df8c",
   134 => x"0c80df88",
   135 => x"08810580",
   136 => x"df880c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"df900cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"df900c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280df",
   177 => x"90088407",
   178 => x"80df900c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80da",
   183 => x"900c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80df90",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80de",
   208 => x"f80c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02f4050d",
  1093 => x"74765452",
  1094 => x"72708105",
  1095 => x"5480f52d",
  1096 => x"51707270",
  1097 => x"81055481",
  1098 => x"b72d70ec",
  1099 => x"38707281",
  1100 => x"b72d028c",
  1101 => x"050d0402",
  1102 => x"f4050d80",
  1103 => x"daac0b80",
  1104 => x"f52d80dd",
  1105 => x"94087081",
  1106 => x"06535452",
  1107 => x"70802e85",
  1108 => x"38718407",
  1109 => x"5272812a",
  1110 => x"70810651",
  1111 => x"5170802e",
  1112 => x"85387182",
  1113 => x"07527282",
  1114 => x"2a708106",
  1115 => x"51517080",
  1116 => x"2e853871",
  1117 => x"81075272",
  1118 => x"832a7081",
  1119 => x"06515170",
  1120 => x"802e8538",
  1121 => x"71880752",
  1122 => x"72842a70",
  1123 => x"81065151",
  1124 => x"70802e85",
  1125 => x"38719007",
  1126 => x"5272852a",
  1127 => x"70810651",
  1128 => x"5170802e",
  1129 => x"853871a0",
  1130 => x"07527288",
  1131 => x"2a708106",
  1132 => x"51517080",
  1133 => x"2e863871",
  1134 => x"80c00752",
  1135 => x"72892a70",
  1136 => x"81065151",
  1137 => x"70802e86",
  1138 => x"38718180",
  1139 => x"075271fc",
  1140 => x"0c7180de",
  1141 => x"f80c028c",
  1142 => x"050d0402",
  1143 => x"cc050d7e",
  1144 => x"5d800b80",
  1145 => x"dd940881",
  1146 => x"8006715c",
  1147 => x"5d5b810b",
  1148 => x"ec0c840b",
  1149 => x"ec0c7c52",
  1150 => x"80df9451",
  1151 => x"80ccad2d",
  1152 => x"80def808",
  1153 => x"7b2e80ff",
  1154 => x"3880df98",
  1155 => x"087bff12",
  1156 => x"57595774",
  1157 => x"7b2e8b38",
  1158 => x"81187581",
  1159 => x"2a565874",
  1160 => x"f738f718",
  1161 => x"58815b80",
  1162 => x"772580db",
  1163 => x"38775274",
  1164 => x"5184a82d",
  1165 => x"80dfe852",
  1166 => x"80df9451",
  1167 => x"80cf822d",
  1168 => x"80def808",
  1169 => x"802ea638",
  1170 => x"80dfe859",
  1171 => x"7ba73883",
  1172 => x"ff567870",
  1173 => x"81055a80",
  1174 => x"f52d7a81",
  1175 => x"1c5ce40c",
  1176 => x"e80cff16",
  1177 => x"56758025",
  1178 => x"e938a4f5",
  1179 => x"0480def8",
  1180 => x"085b8480",
  1181 => x"5780df94",
  1182 => x"5180ced1",
  1183 => x"2dfc8017",
  1184 => x"81165657",
  1185 => x"a4a70480",
  1186 => x"df9808f8",
  1187 => x"0c881d54",
  1188 => x"807480f5",
  1189 => x"2d7081ff",
  1190 => x"06555855",
  1191 => x"72752eb6",
  1192 => x"38811480",
  1193 => x"f52d5372",
  1194 => x"752eab38",
  1195 => x"74821580",
  1196 => x"f52d5456",
  1197 => x"7280d32e",
  1198 => x"09810683",
  1199 => x"38815672",
  1200 => x"80f33270",
  1201 => x"09810570",
  1202 => x"80257807",
  1203 => x"51515372",
  1204 => x"802e8338",
  1205 => x"a0558077",
  1206 => x"81ff0654",
  1207 => x"567280c5",
  1208 => x"2e098106",
  1209 => x"83388156",
  1210 => x"7280e532",
  1211 => x"70098105",
  1212 => x"70802578",
  1213 => x"07515153",
  1214 => x"72802ea4",
  1215 => x"38811480",
  1216 => x"f52d5372",
  1217 => x"b02e0981",
  1218 => x"06893874",
  1219 => x"82800755",
  1220 => x"a6a00472",
  1221 => x"b72e0981",
  1222 => x"06863874",
  1223 => x"84800755",
  1224 => x"80dd9408",
  1225 => x"f9df0675",
  1226 => x"0780dd94",
  1227 => x"0ca2b72d",
  1228 => x"800be00c",
  1229 => x"805186da",
  1230 => x"2d86c72d",
  1231 => x"7a802e88",
  1232 => x"3880da98",
  1233 => x"51a6cc04",
  1234 => x"80dbc051",
  1235 => x"b0d42d7a",
  1236 => x"80def80c",
  1237 => x"02b4050d",
  1238 => x"0402f405",
  1239 => x"0d840bec",
  1240 => x"0c810be0",
  1241 => x"0cae912d",
  1242 => x"a7eb2d81",
  1243 => x"f92d8352",
  1244 => x"adf42d81",
  1245 => x"51858d2d",
  1246 => x"ff125271",
  1247 => x"8025f138",
  1248 => x"840bec0c",
  1249 => x"80d8bc51",
  1250 => x"86a02d80",
  1251 => x"c2d22d80",
  1252 => x"def80880",
  1253 => x"2ebe38a3",
  1254 => x"db5180d6",
  1255 => x"dd2d80da",
  1256 => x"9851b0d4",
  1257 => x"2daeb32d",
  1258 => x"a9962d80",
  1259 => x"def80881",
  1260 => x"06527180",
  1261 => x"2e863880",
  1262 => x"5194bf2d",
  1263 => x"b0e72d80",
  1264 => x"def80852",
  1265 => x"a2b72d86",
  1266 => x"53718338",
  1267 => x"845372ec",
  1268 => x"0ca7a804",
  1269 => x"800b80de",
  1270 => x"f80c028c",
  1271 => x"050d0471",
  1272 => x"980c04ff",
  1273 => x"b00880de",
  1274 => x"f80c0481",
  1275 => x"0bffb00c",
  1276 => x"04800bff",
  1277 => x"b00c0402",
  1278 => x"d8050dff",
  1279 => x"b40887ff",
  1280 => x"ff065a81",
  1281 => x"54807080",
  1282 => x"dd800880",
  1283 => x"dd840880",
  1284 => x"dcdc5b59",
  1285 => x"575a5879",
  1286 => x"74067575",
  1287 => x"06525271",
  1288 => x"712e8d38",
  1289 => x"8077818a",
  1290 => x"2d730975",
  1291 => x"06720755",
  1292 => x"7680e02d",
  1293 => x"7083ffff",
  1294 => x"06535171",
  1295 => x"80e42e09",
  1296 => x"8106a238",
  1297 => x"74740670",
  1298 => x"77760632",
  1299 => x"70098105",
  1300 => x"7072079f",
  1301 => x"2a7b0577",
  1302 => x"097a0674",
  1303 => x"075a5b53",
  1304 => x"5353a8f3",
  1305 => x"047180e4",
  1306 => x"26893881",
  1307 => x"11517077",
  1308 => x"818a2d73",
  1309 => x"10811a82",
  1310 => x"19595a54",
  1311 => x"907925ff",
  1312 => x"96387580",
  1313 => x"dd840c74",
  1314 => x"80dd800c",
  1315 => x"7780def8",
  1316 => x"0c02a805",
  1317 => x"0d0402d0",
  1318 => x"050d805c",
  1319 => x"aaa60480",
  1320 => x"def80881",
  1321 => x"f02e0981",
  1322 => x"068a3881",
  1323 => x"0b80dd8c",
  1324 => x"0caaa604",
  1325 => x"80def808",
  1326 => x"81e02e09",
  1327 => x"81068a38",
  1328 => x"810b80dd",
  1329 => x"900caaa6",
  1330 => x"0480def8",
  1331 => x"085280dd",
  1332 => x"9008802e",
  1333 => x"893880de",
  1334 => x"f8088180",
  1335 => x"05527184",
  1336 => x"2c728f06",
  1337 => x"535380dd",
  1338 => x"8c08802e",
  1339 => x"9a387284",
  1340 => x"2980dbe4",
  1341 => x"05721381",
  1342 => x"712b7009",
  1343 => x"73080673",
  1344 => x"0c515353",
  1345 => x"aa9a0472",
  1346 => x"842980db",
  1347 => x"e4057213",
  1348 => x"83712b72",
  1349 => x"0807720c",
  1350 => x"5353800b",
  1351 => x"80dd900c",
  1352 => x"800b80dd",
  1353 => x"8c0c80df",
  1354 => x"a051ace7",
  1355 => x"2d80def8",
  1356 => x"08ff24fe",
  1357 => x"ea38a7f7",
  1358 => x"2d80def8",
  1359 => x"08802e81",
  1360 => x"b0388159",
  1361 => x"800b80dd",
  1362 => x"880880dd",
  1363 => x"840880dc",
  1364 => x"b85a5c5c",
  1365 => x"587a7906",
  1366 => x"7a7a0654",
  1367 => x"5271732e",
  1368 => x"80f83872",
  1369 => x"09810570",
  1370 => x"74078025",
  1371 => x"80dca41a",
  1372 => x"80f52d70",
  1373 => x"842c718f",
  1374 => x"06585357",
  1375 => x"57527580",
  1376 => x"2ea33871",
  1377 => x"842980db",
  1378 => x"e4057415",
  1379 => x"83712b72",
  1380 => x"0807720c",
  1381 => x"54527680",
  1382 => x"e02d8105",
  1383 => x"52717781",
  1384 => x"8a2dabbb",
  1385 => x"04718429",
  1386 => x"80dbe405",
  1387 => x"74158171",
  1388 => x"2b700973",
  1389 => x"0806730c",
  1390 => x"51535374",
  1391 => x"85327009",
  1392 => x"81057080",
  1393 => x"25515152",
  1394 => x"75802e8e",
  1395 => x"38817073",
  1396 => x"06535371",
  1397 => x"802e8338",
  1398 => x"725c7810",
  1399 => x"81198219",
  1400 => x"59595990",
  1401 => x"7825feed",
  1402 => x"3880dd84",
  1403 => x"0880dd88",
  1404 => x"0c7b80de",
  1405 => x"f80c02b0",
  1406 => x"050d0402",
  1407 => x"f8050d80",
  1408 => x"dbe4528f",
  1409 => x"51807270",
  1410 => x"8405540c",
  1411 => x"ff115170",
  1412 => x"8025f238",
  1413 => x"0288050d",
  1414 => x"0402f005",
  1415 => x"0d7551a7",
  1416 => x"f12d7082",
  1417 => x"2cfc0680",
  1418 => x"dbe41172",
  1419 => x"109e0671",
  1420 => x"0870722a",
  1421 => x"70830682",
  1422 => x"742b7009",
  1423 => x"7406760c",
  1424 => x"54515657",
  1425 => x"535153a7",
  1426 => x"eb2d7180",
  1427 => x"def80c02",
  1428 => x"90050d04",
  1429 => x"02fc050d",
  1430 => x"72518071",
  1431 => x"0c800b84",
  1432 => x"120c0284",
  1433 => x"050d0402",
  1434 => x"f0050d75",
  1435 => x"70088412",
  1436 => x"08535353",
  1437 => x"ff547171",
  1438 => x"2ea838a7",
  1439 => x"f12d8413",
  1440 => x"08708429",
  1441 => x"14881170",
  1442 => x"087081ff",
  1443 => x"06841808",
  1444 => x"81118706",
  1445 => x"841a0c53",
  1446 => x"51555151",
  1447 => x"51a7eb2d",
  1448 => x"71547380",
  1449 => x"def80c02",
  1450 => x"90050d04",
  1451 => x"02f8050d",
  1452 => x"a7f12de0",
  1453 => x"08708b2a",
  1454 => x"70810651",
  1455 => x"52527080",
  1456 => x"2ea13880",
  1457 => x"dfa00870",
  1458 => x"842980df",
  1459 => x"a8057381",
  1460 => x"ff06710c",
  1461 => x"515180df",
  1462 => x"a0088111",
  1463 => x"870680df",
  1464 => x"a00c5180",
  1465 => x"0b80dfc8",
  1466 => x"0ca7e32d",
  1467 => x"a7eb2d02",
  1468 => x"88050d04",
  1469 => x"02fc050d",
  1470 => x"a7f12d81",
  1471 => x"0b80dfc8",
  1472 => x"0ca7eb2d",
  1473 => x"80dfc808",
  1474 => x"5170f938",
  1475 => x"0284050d",
  1476 => x"0402fc05",
  1477 => x"0d80dfa0",
  1478 => x"51acd42d",
  1479 => x"abfb2dad",
  1480 => x"ac51a7df",
  1481 => x"2d028405",
  1482 => x"0d0480df",
  1483 => x"d40880de",
  1484 => x"f80c0402",
  1485 => x"fc050d81",
  1486 => x"0b80dd98",
  1487 => x"0c815185",
  1488 => x"8d2d0284",
  1489 => x"050d0402",
  1490 => x"fc050dae",
  1491 => x"d104a996",
  1492 => x"2d80f651",
  1493 => x"ac992d80",
  1494 => x"def808f2",
  1495 => x"3880da51",
  1496 => x"ac992d80",
  1497 => x"def808e6",
  1498 => x"3880def8",
  1499 => x"0880dd98",
  1500 => x"0c80def8",
  1501 => x"0851858d",
  1502 => x"2d028405",
  1503 => x"0d0402ec",
  1504 => x"050d7654",
  1505 => x"8052870b",
  1506 => x"881580f5",
  1507 => x"2d565374",
  1508 => x"72248338",
  1509 => x"a0537251",
  1510 => x"83842d81",
  1511 => x"128b1580",
  1512 => x"f52d5452",
  1513 => x"727225de",
  1514 => x"38029405",
  1515 => x"0d0402f0",
  1516 => x"050d80df",
  1517 => x"d4085481",
  1518 => x"f92d800b",
  1519 => x"80dfd80c",
  1520 => x"7308802e",
  1521 => x"81893882",
  1522 => x"0b80df8c",
  1523 => x"0c80dfd8",
  1524 => x"088f0680",
  1525 => x"df880c73",
  1526 => x"08527183",
  1527 => x"2e963871",
  1528 => x"83268938",
  1529 => x"71812eb0",
  1530 => x"38b0b804",
  1531 => x"71852ea0",
  1532 => x"38b0b804",
  1533 => x"881480f5",
  1534 => x"2d841508",
  1535 => x"80d8d453",
  1536 => x"545286a0",
  1537 => x"2d718429",
  1538 => x"13700852",
  1539 => x"52b0bc04",
  1540 => x"7351aefe",
  1541 => x"2db0b804",
  1542 => x"80dd9408",
  1543 => x"8815082c",
  1544 => x"70810651",
  1545 => x"5271802e",
  1546 => x"883880d8",
  1547 => x"d851b0b5",
  1548 => x"0480d8dc",
  1549 => x"5186a02d",
  1550 => x"84140851",
  1551 => x"86a02d80",
  1552 => x"dfd80881",
  1553 => x"0580dfd8",
  1554 => x"0c8c1454",
  1555 => x"afc00402",
  1556 => x"90050d04",
  1557 => x"7180dfd4",
  1558 => x"0cafae2d",
  1559 => x"80dfd808",
  1560 => x"ff0580df",
  1561 => x"dc0c0402",
  1562 => x"e8050d80",
  1563 => x"dfd40880",
  1564 => x"dfe00857",
  1565 => x"5580f651",
  1566 => x"ac992d80",
  1567 => x"def80881",
  1568 => x"2a708106",
  1569 => x"51527180",
  1570 => x"2ea438b1",
  1571 => x"9104a996",
  1572 => x"2d80f651",
  1573 => x"ac992d80",
  1574 => x"def808f2",
  1575 => x"3880dd98",
  1576 => x"08813270",
  1577 => x"80dd980c",
  1578 => x"70525285",
  1579 => x"8d2d800b",
  1580 => x"80dfcc0c",
  1581 => x"800b80df",
  1582 => x"d00c80dd",
  1583 => x"9808838d",
  1584 => x"3880da51",
  1585 => x"ac992d80",
  1586 => x"def80880",
  1587 => x"2e8c3880",
  1588 => x"dfcc0881",
  1589 => x"800780df",
  1590 => x"cc0c80d9",
  1591 => x"51ac992d",
  1592 => x"80def808",
  1593 => x"802e8c38",
  1594 => x"80dfcc08",
  1595 => x"80c00780",
  1596 => x"dfcc0c81",
  1597 => x"9451ac99",
  1598 => x"2d80def8",
  1599 => x"08802e8b",
  1600 => x"3880dfcc",
  1601 => x"08900780",
  1602 => x"dfcc0c81",
  1603 => x"9151ac99",
  1604 => x"2d80def8",
  1605 => x"08802e8b",
  1606 => x"3880dfcc",
  1607 => x"08a00780",
  1608 => x"dfcc0c81",
  1609 => x"f551ac99",
  1610 => x"2d80def8",
  1611 => x"08802e8b",
  1612 => x"3880dfcc",
  1613 => x"08810780",
  1614 => x"dfcc0c81",
  1615 => x"f251ac99",
  1616 => x"2d80def8",
  1617 => x"08802e8b",
  1618 => x"3880dfcc",
  1619 => x"08820780",
  1620 => x"dfcc0c81",
  1621 => x"eb51ac99",
  1622 => x"2d80def8",
  1623 => x"08802e8b",
  1624 => x"3880dfcc",
  1625 => x"08840780",
  1626 => x"dfcc0c81",
  1627 => x"f451ac99",
  1628 => x"2d80def8",
  1629 => x"08802e8b",
  1630 => x"3880dfcc",
  1631 => x"08880780",
  1632 => x"dfcc0c80",
  1633 => x"d851ac99",
  1634 => x"2d80def8",
  1635 => x"08802e8c",
  1636 => x"3880dfd0",
  1637 => x"08818007",
  1638 => x"80dfd00c",
  1639 => x"9251ac99",
  1640 => x"2d80def8",
  1641 => x"08802e8c",
  1642 => x"3880dfd0",
  1643 => x"0880c007",
  1644 => x"80dfd00c",
  1645 => x"9451ac99",
  1646 => x"2d80def8",
  1647 => x"08802e8b",
  1648 => x"3880dfd0",
  1649 => x"08900780",
  1650 => x"dfd00c91",
  1651 => x"51ac992d",
  1652 => x"80def808",
  1653 => x"802e8b38",
  1654 => x"80dfd008",
  1655 => x"a00780df",
  1656 => x"d00c9d51",
  1657 => x"ac992d80",
  1658 => x"def80880",
  1659 => x"2e8b3880",
  1660 => x"dfd00881",
  1661 => x"0780dfd0",
  1662 => x"0c9b51ac",
  1663 => x"992d80de",
  1664 => x"f808802e",
  1665 => x"8b3880df",
  1666 => x"d0088207",
  1667 => x"80dfd00c",
  1668 => x"9c51ac99",
  1669 => x"2d80def8",
  1670 => x"08802e8b",
  1671 => x"3880dfd0",
  1672 => x"08840780",
  1673 => x"dfd00ca3",
  1674 => x"51ac992d",
  1675 => x"80def808",
  1676 => x"802e8b38",
  1677 => x"80dfd008",
  1678 => x"880780df",
  1679 => x"d00c81fd",
  1680 => x"51ac992d",
  1681 => x"81fa51ac",
  1682 => x"992dbaa2",
  1683 => x"0481f551",
  1684 => x"ac992d80",
  1685 => x"def80881",
  1686 => x"2a708106",
  1687 => x"51527180",
  1688 => x"2eb33880",
  1689 => x"dfdc0852",
  1690 => x"71802e8a",
  1691 => x"38ff1280",
  1692 => x"dfdc0cb5",
  1693 => x"950480df",
  1694 => x"d8081080",
  1695 => x"dfd80805",
  1696 => x"70842916",
  1697 => x"51528812",
  1698 => x"08802e89",
  1699 => x"38ff5188",
  1700 => x"12085271",
  1701 => x"2d81f251",
  1702 => x"ac992d80",
  1703 => x"def80881",
  1704 => x"2a708106",
  1705 => x"51527180",
  1706 => x"2eb43880",
  1707 => x"dfd808ff",
  1708 => x"1180dfdc",
  1709 => x"08565353",
  1710 => x"7372258a",
  1711 => x"38811480",
  1712 => x"dfdc0cb5",
  1713 => x"de047210",
  1714 => x"13708429",
  1715 => x"16515288",
  1716 => x"1208802e",
  1717 => x"8938fe51",
  1718 => x"88120852",
  1719 => x"712d81fd",
  1720 => x"51ac992d",
  1721 => x"80def808",
  1722 => x"812a7081",
  1723 => x"06515271",
  1724 => x"802eb138",
  1725 => x"80dfdc08",
  1726 => x"802e8a38",
  1727 => x"800b80df",
  1728 => x"dc0cb6a4",
  1729 => x"0480dfd8",
  1730 => x"081080df",
  1731 => x"d8080570",
  1732 => x"84291651",
  1733 => x"52881208",
  1734 => x"802e8938",
  1735 => x"fd518812",
  1736 => x"0852712d",
  1737 => x"81fa51ac",
  1738 => x"992d80de",
  1739 => x"f808812a",
  1740 => x"70810651",
  1741 => x"5271802e",
  1742 => x"b13880df",
  1743 => x"d808ff11",
  1744 => x"545280df",
  1745 => x"dc087325",
  1746 => x"89387280",
  1747 => x"dfdc0cb6",
  1748 => x"ea047110",
  1749 => x"12708429",
  1750 => x"16515288",
  1751 => x"1208802e",
  1752 => x"8938fc51",
  1753 => x"88120852",
  1754 => x"712d80df",
  1755 => x"dc087053",
  1756 => x"5473802e",
  1757 => x"8a388c15",
  1758 => x"ff155555",
  1759 => x"b6f10482",
  1760 => x"0b80df8c",
  1761 => x"0c718f06",
  1762 => x"80df880c",
  1763 => x"81eb51ac",
  1764 => x"992d80de",
  1765 => x"f808812a",
  1766 => x"70810651",
  1767 => x"5271802e",
  1768 => x"ad387408",
  1769 => x"852e0981",
  1770 => x"06a43888",
  1771 => x"1580f52d",
  1772 => x"ff055271",
  1773 => x"881681b7",
  1774 => x"2d71982b",
  1775 => x"52718025",
  1776 => x"8838800b",
  1777 => x"881681b7",
  1778 => x"2d7451ae",
  1779 => x"fe2d81f4",
  1780 => x"51ac992d",
  1781 => x"80def808",
  1782 => x"812a7081",
  1783 => x"06515271",
  1784 => x"802eb338",
  1785 => x"7408852e",
  1786 => x"098106aa",
  1787 => x"38881580",
  1788 => x"f52d8105",
  1789 => x"52718816",
  1790 => x"81b72d71",
  1791 => x"81ff068b",
  1792 => x"1680f52d",
  1793 => x"54527272",
  1794 => x"27873872",
  1795 => x"881681b7",
  1796 => x"2d7451ae",
  1797 => x"fe2d80da",
  1798 => x"51ac992d",
  1799 => x"80def808",
  1800 => x"812a7081",
  1801 => x"06515271",
  1802 => x"802e81ad",
  1803 => x"3880dfd4",
  1804 => x"0880dfdc",
  1805 => x"08555373",
  1806 => x"802e8a38",
  1807 => x"8c13ff15",
  1808 => x"5553b8b7",
  1809 => x"04720852",
  1810 => x"71822ea6",
  1811 => x"38718226",
  1812 => x"89387181",
  1813 => x"2eaa38b9",
  1814 => x"d9047183",
  1815 => x"2eb43871",
  1816 => x"842e0981",
  1817 => x"0680f238",
  1818 => x"88130851",
  1819 => x"b0d42db9",
  1820 => x"d90480df",
  1821 => x"dc085188",
  1822 => x"13085271",
  1823 => x"2db9d904",
  1824 => x"810b8814",
  1825 => x"082b80dd",
  1826 => x"94083280",
  1827 => x"dd940cb9",
  1828 => x"ad048813",
  1829 => x"80f52d81",
  1830 => x"058b1480",
  1831 => x"f52d5354",
  1832 => x"71742483",
  1833 => x"38805473",
  1834 => x"881481b7",
  1835 => x"2dafae2d",
  1836 => x"b9d90475",
  1837 => x"08802ea4",
  1838 => x"38750851",
  1839 => x"ac992d80",
  1840 => x"def80881",
  1841 => x"06527180",
  1842 => x"2e8c3880",
  1843 => x"dfdc0851",
  1844 => x"84160852",
  1845 => x"712d8816",
  1846 => x"5675d838",
  1847 => x"8054800b",
  1848 => x"80df8c0c",
  1849 => x"738f0680",
  1850 => x"df880ca0",
  1851 => x"527380df",
  1852 => x"dc082e09",
  1853 => x"81069938",
  1854 => x"80dfd808",
  1855 => x"ff057432",
  1856 => x"70098105",
  1857 => x"7072079f",
  1858 => x"2a917131",
  1859 => x"51515353",
  1860 => x"71518384",
  1861 => x"2d811454",
  1862 => x"8e7425c2",
  1863 => x"3880dd98",
  1864 => x"08527180",
  1865 => x"def80c02",
  1866 => x"98050d04",
  1867 => x"02f4050d",
  1868 => x"d45281ff",
  1869 => x"720c7108",
  1870 => x"5381ff72",
  1871 => x"0c72882b",
  1872 => x"83fe8006",
  1873 => x"72087081",
  1874 => x"ff065152",
  1875 => x"5381ff72",
  1876 => x"0c727107",
  1877 => x"882b7208",
  1878 => x"7081ff06",
  1879 => x"51525381",
  1880 => x"ff720c72",
  1881 => x"7107882b",
  1882 => x"72087081",
  1883 => x"ff067207",
  1884 => x"80def80c",
  1885 => x"5253028c",
  1886 => x"050d0402",
  1887 => x"f4050d74",
  1888 => x"767181ff",
  1889 => x"06d40c53",
  1890 => x"5380dfe4",
  1891 => x"08853871",
  1892 => x"892b5271",
  1893 => x"982ad40c",
  1894 => x"71902a70",
  1895 => x"81ff06d4",
  1896 => x"0c517188",
  1897 => x"2a7081ff",
  1898 => x"06d40c51",
  1899 => x"7181ff06",
  1900 => x"d40c7290",
  1901 => x"2a7081ff",
  1902 => x"06d40c51",
  1903 => x"d4087081",
  1904 => x"ff065151",
  1905 => x"82b8bf52",
  1906 => x"7081ff2e",
  1907 => x"09810694",
  1908 => x"3881ff0b",
  1909 => x"d40cd408",
  1910 => x"7081ff06",
  1911 => x"ff145451",
  1912 => x"5171e538",
  1913 => x"7080def8",
  1914 => x"0c028c05",
  1915 => x"0d0402fc",
  1916 => x"050d81c7",
  1917 => x"5181ff0b",
  1918 => x"d40cff11",
  1919 => x"51708025",
  1920 => x"f4380284",
  1921 => x"050d0402",
  1922 => x"f4050d81",
  1923 => x"ff0bd40c",
  1924 => x"93538052",
  1925 => x"87fc80c1",
  1926 => x"51bafb2d",
  1927 => x"80def808",
  1928 => x"8b3881ff",
  1929 => x"0bd40c81",
  1930 => x"53bcb504",
  1931 => x"bbee2dff",
  1932 => x"135372de",
  1933 => x"387280de",
  1934 => x"f80c028c",
  1935 => x"050d0402",
  1936 => x"ec050d81",
  1937 => x"0b80dfe4",
  1938 => x"0c8454d0",
  1939 => x"08708f2a",
  1940 => x"70810651",
  1941 => x"515372f3",
  1942 => x"3872d00c",
  1943 => x"bbee2d80",
  1944 => x"d8e05186",
  1945 => x"a02dd008",
  1946 => x"708f2a70",
  1947 => x"81065151",
  1948 => x"5372f338",
  1949 => x"810bd00c",
  1950 => x"b1538052",
  1951 => x"84d480c0",
  1952 => x"51bafb2d",
  1953 => x"80def808",
  1954 => x"812e9338",
  1955 => x"72822ebf",
  1956 => x"38ff1353",
  1957 => x"72e438ff",
  1958 => x"145473ff",
  1959 => x"ae38bbee",
  1960 => x"2d83aa52",
  1961 => x"849c80c8",
  1962 => x"51bafb2d",
  1963 => x"80def808",
  1964 => x"812e0981",
  1965 => x"069338ba",
  1966 => x"ac2d80de",
  1967 => x"f80883ff",
  1968 => x"ff065372",
  1969 => x"83aa2e9f",
  1970 => x"38bc872d",
  1971 => x"bde20480",
  1972 => x"d8ec5186",
  1973 => x"a02d8053",
  1974 => x"bfb70480",
  1975 => x"d9845186",
  1976 => x"a02d8054",
  1977 => x"bf880481",
  1978 => x"ff0bd40c",
  1979 => x"b154bbee",
  1980 => x"2d8fcf53",
  1981 => x"805287fc",
  1982 => x"80f751ba",
  1983 => x"fb2d80de",
  1984 => x"f8085580",
  1985 => x"def80881",
  1986 => x"2e098106",
  1987 => x"9c3881ff",
  1988 => x"0bd40c82",
  1989 => x"0a52849c",
  1990 => x"80e951ba",
  1991 => x"fb2d80de",
  1992 => x"f808802e",
  1993 => x"8d38bbee",
  1994 => x"2dff1353",
  1995 => x"72c638be",
  1996 => x"fb0481ff",
  1997 => x"0bd40c80",
  1998 => x"def80852",
  1999 => x"87fc80fa",
  2000 => x"51bafb2d",
  2001 => x"80def808",
  2002 => x"b23881ff",
  2003 => x"0bd40cd4",
  2004 => x"085381ff",
  2005 => x"0bd40c81",
  2006 => x"ff0bd40c",
  2007 => x"81ff0bd4",
  2008 => x"0c81ff0b",
  2009 => x"d40c7286",
  2010 => x"2a708106",
  2011 => x"76565153",
  2012 => x"72963880",
  2013 => x"def80854",
  2014 => x"bf880473",
  2015 => x"822efedb",
  2016 => x"38ff1454",
  2017 => x"73fee738",
  2018 => x"7380dfe4",
  2019 => x"0c738b38",
  2020 => x"815287fc",
  2021 => x"80d051ba",
  2022 => x"fb2d81ff",
  2023 => x"0bd40cd0",
  2024 => x"08708f2a",
  2025 => x"70810651",
  2026 => x"515372f3",
  2027 => x"3872d00c",
  2028 => x"81ff0bd4",
  2029 => x"0c815372",
  2030 => x"80def80c",
  2031 => x"0294050d",
  2032 => x"0402e805",
  2033 => x"0d785580",
  2034 => x"5681ff0b",
  2035 => x"d40cd008",
  2036 => x"708f2a70",
  2037 => x"81065151",
  2038 => x"5372f338",
  2039 => x"82810bd0",
  2040 => x"0c81ff0b",
  2041 => x"d40c7752",
  2042 => x"87fc80d1",
  2043 => x"51bafb2d",
  2044 => x"80dbc6df",
  2045 => x"5480def8",
  2046 => x"08802e8c",
  2047 => x"3880d9a4",
  2048 => x"5186a02d",
  2049 => x"80c0dd04",
  2050 => x"81ff0bd4",
  2051 => x"0cd40870",
  2052 => x"81ff0651",
  2053 => x"537281fe",
  2054 => x"2e098106",
  2055 => x"9f3880ff",
  2056 => x"53baac2d",
  2057 => x"80def808",
  2058 => x"75708405",
  2059 => x"570cff13",
  2060 => x"53728025",
  2061 => x"ec388156",
  2062 => x"80c0c204",
  2063 => x"ff145473",
  2064 => x"c73881ff",
  2065 => x"0bd40c81",
  2066 => x"ff0bd40c",
  2067 => x"d008708f",
  2068 => x"2a708106",
  2069 => x"51515372",
  2070 => x"f33872d0",
  2071 => x"0c7580de",
  2072 => x"f80c0298",
  2073 => x"050d0402",
  2074 => x"e8050d77",
  2075 => x"797b5855",
  2076 => x"55805372",
  2077 => x"7625a538",
  2078 => x"74708105",
  2079 => x"5680f52d",
  2080 => x"74708105",
  2081 => x"5680f52d",
  2082 => x"52527171",
  2083 => x"2e873881",
  2084 => x"5180c19e",
  2085 => x"04811353",
  2086 => x"80c0f304",
  2087 => x"80517080",
  2088 => x"def80c02",
  2089 => x"98050d04",
  2090 => x"02ec050d",
  2091 => x"76557480",
  2092 => x"2e80c438",
  2093 => x"9a1580e0",
  2094 => x"2d5180cf",
  2095 => x"dc2d80de",
  2096 => x"f80880de",
  2097 => x"f80880e6",
  2098 => x"980c80de",
  2099 => x"f8085454",
  2100 => x"80e5f408",
  2101 => x"802e9b38",
  2102 => x"941580e0",
  2103 => x"2d5180cf",
  2104 => x"dc2d80de",
  2105 => x"f808902b",
  2106 => x"83fff00a",
  2107 => x"06707507",
  2108 => x"51537280",
  2109 => x"e6980c80",
  2110 => x"e6980853",
  2111 => x"72802e9e",
  2112 => x"3880e5ec",
  2113 => x"08fe1471",
  2114 => x"2980e680",
  2115 => x"080580e6",
  2116 => x"9c0c7084",
  2117 => x"2b80e5f8",
  2118 => x"0c5480c2",
  2119 => x"cd0480e6",
  2120 => x"840880e6",
  2121 => x"980c80e6",
  2122 => x"880880e6",
  2123 => x"9c0c80e5",
  2124 => x"f408802e",
  2125 => x"8c3880e5",
  2126 => x"ec08842b",
  2127 => x"5380c2c8",
  2128 => x"0480e68c",
  2129 => x"08842b53",
  2130 => x"7280e5f8",
  2131 => x"0c029405",
  2132 => x"0d0402d8",
  2133 => x"050d800b",
  2134 => x"80e5f40c",
  2135 => x"8454bcbf",
  2136 => x"2d80def8",
  2137 => x"08802e98",
  2138 => x"3880dfe8",
  2139 => x"528051bf",
  2140 => x"c12d80de",
  2141 => x"f808802e",
  2142 => x"8738fe54",
  2143 => x"80c38804",
  2144 => x"ff145473",
  2145 => x"8024d738",
  2146 => x"738e3880",
  2147 => x"d9b45186",
  2148 => x"a02d7355",
  2149 => x"80c8eb04",
  2150 => x"8056810b",
  2151 => x"80e6a00c",
  2152 => x"885380d9",
  2153 => x"c85280e0",
  2154 => x"9e5180c0",
  2155 => x"e72d80de",
  2156 => x"f808762e",
  2157 => x"09810689",
  2158 => x"3880def8",
  2159 => x"0880e6a0",
  2160 => x"0c885380",
  2161 => x"d9d45280",
  2162 => x"e0ba5180",
  2163 => x"c0e72d80",
  2164 => x"def80889",
  2165 => x"3880def8",
  2166 => x"0880e6a0",
  2167 => x"0c80e6a0",
  2168 => x"08802e81",
  2169 => x"843880e3",
  2170 => x"ae0b80f5",
  2171 => x"2d80e3af",
  2172 => x"0b80f52d",
  2173 => x"71982b71",
  2174 => x"902b0780",
  2175 => x"e3b00b80",
  2176 => x"f52d7088",
  2177 => x"2b720780",
  2178 => x"e3b10b80",
  2179 => x"f52d7107",
  2180 => x"80e3e60b",
  2181 => x"80f52d80",
  2182 => x"e3e70b80",
  2183 => x"f52d7188",
  2184 => x"2b07535f",
  2185 => x"54525a56",
  2186 => x"57557381",
  2187 => x"abaa2e09",
  2188 => x"81069038",
  2189 => x"755180cf",
  2190 => x"ab2d80de",
  2191 => x"f8085680",
  2192 => x"c4d20473",
  2193 => x"82d4d52e",
  2194 => x"893880d9",
  2195 => x"e05180c5",
  2196 => x"a10480df",
  2197 => x"e8527551",
  2198 => x"bfc12d80",
  2199 => x"def80855",
  2200 => x"80def808",
  2201 => x"802e8483",
  2202 => x"38885380",
  2203 => x"d9d45280",
  2204 => x"e0ba5180",
  2205 => x"c0e72d80",
  2206 => x"def8088b",
  2207 => x"38810b80",
  2208 => x"e5f40c80",
  2209 => x"c5a80488",
  2210 => x"5380d9c8",
  2211 => x"5280e09e",
  2212 => x"5180c0e7",
  2213 => x"2d80def8",
  2214 => x"08802e8c",
  2215 => x"3880d9f4",
  2216 => x"5186a02d",
  2217 => x"80c68704",
  2218 => x"80e3e60b",
  2219 => x"80f52d54",
  2220 => x"7380d52e",
  2221 => x"09810680",
  2222 => x"ce3880e3",
  2223 => x"e70b80f5",
  2224 => x"2d547381",
  2225 => x"aa2e0981",
  2226 => x"06bd3880",
  2227 => x"0b80dfe8",
  2228 => x"0b80f52d",
  2229 => x"56547481",
  2230 => x"e92e8338",
  2231 => x"81547481",
  2232 => x"eb2e8c38",
  2233 => x"80557375",
  2234 => x"2e098106",
  2235 => x"82fd3880",
  2236 => x"dff30b80",
  2237 => x"f52d5574",
  2238 => x"8e3880df",
  2239 => x"f40b80f5",
  2240 => x"2d547382",
  2241 => x"2e873880",
  2242 => x"5580c8eb",
  2243 => x"0480dff5",
  2244 => x"0b80f52d",
  2245 => x"7080e5ec",
  2246 => x"0cff0580",
  2247 => x"e5f00c80",
  2248 => x"dff60b80",
  2249 => x"f52d80df",
  2250 => x"f70b80f5",
  2251 => x"2d587605",
  2252 => x"77828029",
  2253 => x"057080e5",
  2254 => x"fc0c80df",
  2255 => x"f80b80f5",
  2256 => x"2d7080e6",
  2257 => x"900c80e5",
  2258 => x"f4085957",
  2259 => x"5876802e",
  2260 => x"81b93888",
  2261 => x"5380d9d4",
  2262 => x"5280e0ba",
  2263 => x"5180c0e7",
  2264 => x"2d80def8",
  2265 => x"08828438",
  2266 => x"80e5ec08",
  2267 => x"70842b80",
  2268 => x"e5f80c70",
  2269 => x"80e68c0c",
  2270 => x"80e08d0b",
  2271 => x"80f52d80",
  2272 => x"e08c0b80",
  2273 => x"f52d7182",
  2274 => x"80290580",
  2275 => x"e08e0b80",
  2276 => x"f52d7084",
  2277 => x"80802912",
  2278 => x"80e08f0b",
  2279 => x"80f52d70",
  2280 => x"81800a29",
  2281 => x"127080e6",
  2282 => x"940c80e6",
  2283 => x"90087129",
  2284 => x"80e5fc08",
  2285 => x"057080e6",
  2286 => x"800c80e0",
  2287 => x"950b80f5",
  2288 => x"2d80e094",
  2289 => x"0b80f52d",
  2290 => x"71828029",
  2291 => x"0580e096",
  2292 => x"0b80f52d",
  2293 => x"70848080",
  2294 => x"291280e0",
  2295 => x"970b80f5",
  2296 => x"2d70982b",
  2297 => x"81f00a06",
  2298 => x"72057080",
  2299 => x"e6840cfe",
  2300 => x"117e2977",
  2301 => x"0580e688",
  2302 => x"0c525952",
  2303 => x"43545e51",
  2304 => x"5259525d",
  2305 => x"57595780",
  2306 => x"c8e30480",
  2307 => x"dffa0b80",
  2308 => x"f52d80df",
  2309 => x"f90b80f5",
  2310 => x"2d718280",
  2311 => x"29057080",
  2312 => x"e5f80c70",
  2313 => x"a02983ff",
  2314 => x"0570892a",
  2315 => x"7080e68c",
  2316 => x"0c80dfff",
  2317 => x"0b80f52d",
  2318 => x"80dffe0b",
  2319 => x"80f52d71",
  2320 => x"82802905",
  2321 => x"7080e694",
  2322 => x"0c7b7129",
  2323 => x"1e7080e6",
  2324 => x"880c7d80",
  2325 => x"e6840c73",
  2326 => x"0580e680",
  2327 => x"0c555e51",
  2328 => x"51555580",
  2329 => x"5180c1a8",
  2330 => x"2d815574",
  2331 => x"80def80c",
  2332 => x"02a8050d",
  2333 => x"0402ec05",
  2334 => x"0d767087",
  2335 => x"2c7180ff",
  2336 => x"06555654",
  2337 => x"80e5f408",
  2338 => x"8a387388",
  2339 => x"2c7481ff",
  2340 => x"06545580",
  2341 => x"dfe85280",
  2342 => x"e5fc0815",
  2343 => x"51bfc12d",
  2344 => x"80def808",
  2345 => x"5480def8",
  2346 => x"08802ebb",
  2347 => x"3880e5f4",
  2348 => x"08802e9c",
  2349 => x"38728429",
  2350 => x"80dfe805",
  2351 => x"70085253",
  2352 => x"80cfab2d",
  2353 => x"80def808",
  2354 => x"f00a0653",
  2355 => x"80c9e504",
  2356 => x"721080df",
  2357 => x"e8057080",
  2358 => x"e02d5253",
  2359 => x"80cfdc2d",
  2360 => x"80def808",
  2361 => x"53725473",
  2362 => x"80def80c",
  2363 => x"0294050d",
  2364 => x"0402e005",
  2365 => x"0d797084",
  2366 => x"2c80e69c",
  2367 => x"0805718f",
  2368 => x"06525553",
  2369 => x"728a3880",
  2370 => x"dfe85273",
  2371 => x"51bfc12d",
  2372 => x"72a02980",
  2373 => x"dfe80554",
  2374 => x"807480f5",
  2375 => x"2d565374",
  2376 => x"732e8338",
  2377 => x"81537481",
  2378 => x"e52e81f5",
  2379 => x"38817074",
  2380 => x"06545872",
  2381 => x"802e81e9",
  2382 => x"388b1480",
  2383 => x"f52d7083",
  2384 => x"2a790658",
  2385 => x"56769c38",
  2386 => x"80dd9c08",
  2387 => x"53728938",
  2388 => x"7280e3e8",
  2389 => x"0b81b72d",
  2390 => x"7680dd9c",
  2391 => x"0c735380",
  2392 => x"cca30475",
  2393 => x"8f2e0981",
  2394 => x"0681b638",
  2395 => x"749f068d",
  2396 => x"2980e3db",
  2397 => x"11515381",
  2398 => x"1480f52d",
  2399 => x"73708105",
  2400 => x"5581b72d",
  2401 => x"831480f5",
  2402 => x"2d737081",
  2403 => x"055581b7",
  2404 => x"2d851480",
  2405 => x"f52d7370",
  2406 => x"81055581",
  2407 => x"b72d8714",
  2408 => x"80f52d73",
  2409 => x"70810555",
  2410 => x"81b72d89",
  2411 => x"1480f52d",
  2412 => x"73708105",
  2413 => x"5581b72d",
  2414 => x"8e1480f5",
  2415 => x"2d737081",
  2416 => x"055581b7",
  2417 => x"2d901480",
  2418 => x"f52d7370",
  2419 => x"81055581",
  2420 => x"b72d9214",
  2421 => x"80f52d73",
  2422 => x"70810555",
  2423 => x"81b72d94",
  2424 => x"1480f52d",
  2425 => x"73708105",
  2426 => x"5581b72d",
  2427 => x"961480f5",
  2428 => x"2d737081",
  2429 => x"055581b7",
  2430 => x"2d981480",
  2431 => x"f52d7370",
  2432 => x"81055581",
  2433 => x"b72d9c14",
  2434 => x"80f52d73",
  2435 => x"70810555",
  2436 => x"81b72d9e",
  2437 => x"1480f52d",
  2438 => x"7381b72d",
  2439 => x"7780dd9c",
  2440 => x"0c805372",
  2441 => x"80def80c",
  2442 => x"02a0050d",
  2443 => x"0402cc05",
  2444 => x"0d7e605e",
  2445 => x"5a800b80",
  2446 => x"e6980880",
  2447 => x"e69c0859",
  2448 => x"5c568058",
  2449 => x"80e5f808",
  2450 => x"782e81bd",
  2451 => x"38778f06",
  2452 => x"a0175754",
  2453 => x"73913880",
  2454 => x"dfe85276",
  2455 => x"51811757",
  2456 => x"bfc12d80",
  2457 => x"dfe85680",
  2458 => x"7680f52d",
  2459 => x"56547474",
  2460 => x"2e833881",
  2461 => x"547481e5",
  2462 => x"2e818238",
  2463 => x"81707506",
  2464 => x"555c7380",
  2465 => x"2e80f638",
  2466 => x"8b1680f5",
  2467 => x"2d980659",
  2468 => x"7880ea38",
  2469 => x"8b537c52",
  2470 => x"755180c0",
  2471 => x"e72d80de",
  2472 => x"f80880d9",
  2473 => x"389c1608",
  2474 => x"5180cfab",
  2475 => x"2d80def8",
  2476 => x"08841b0c",
  2477 => x"9a1680e0",
  2478 => x"2d5180cf",
  2479 => x"dc2d80de",
  2480 => x"f80880de",
  2481 => x"f808881c",
  2482 => x"0c80def8",
  2483 => x"08555580",
  2484 => x"e5f40880",
  2485 => x"2e9a3894",
  2486 => x"1680e02d",
  2487 => x"5180cfdc",
  2488 => x"2d80def8",
  2489 => x"08902b83",
  2490 => x"fff00a06",
  2491 => x"70165154",
  2492 => x"73881b0c",
  2493 => x"787a0c7b",
  2494 => x"5480cec7",
  2495 => x"04811858",
  2496 => x"80e5f808",
  2497 => x"7826fec5",
  2498 => x"3880e5f4",
  2499 => x"08802eb5",
  2500 => x"387a5180",
  2501 => x"c8f52d80",
  2502 => x"def80880",
  2503 => x"def80880",
  2504 => x"fffffff8",
  2505 => x"06555b73",
  2506 => x"80ffffff",
  2507 => x"f82e9638",
  2508 => x"80def808",
  2509 => x"fe0580e5",
  2510 => x"ec082980",
  2511 => x"e6800805",
  2512 => x"5780ccc2",
  2513 => x"04805473",
  2514 => x"80def80c",
  2515 => x"02b4050d",
  2516 => x"0402f405",
  2517 => x"0d747008",
  2518 => x"8105710c",
  2519 => x"700880e5",
  2520 => x"f0080653",
  2521 => x"53719038",
  2522 => x"88130851",
  2523 => x"80c8f52d",
  2524 => x"80def808",
  2525 => x"88140c81",
  2526 => x"0b80def8",
  2527 => x"0c028c05",
  2528 => x"0d0402f0",
  2529 => x"050d7588",
  2530 => x"1108fe05",
  2531 => x"80e5ec08",
  2532 => x"2980e680",
  2533 => x"08117208",
  2534 => x"80e5f008",
  2535 => x"06057955",
  2536 => x"535454bf",
  2537 => x"c12d0290",
  2538 => x"050d0402",
  2539 => x"f4050d74",
  2540 => x"70882a83",
  2541 => x"fe800670",
  2542 => x"72982a07",
  2543 => x"72882b87",
  2544 => x"fc808006",
  2545 => x"73982b81",
  2546 => x"f00a0671",
  2547 => x"73070780",
  2548 => x"def80c56",
  2549 => x"51535102",
  2550 => x"8c050d04",
  2551 => x"02f8050d",
  2552 => x"028e0580",
  2553 => x"f52d7488",
  2554 => x"2b077083",
  2555 => x"ffff0680",
  2556 => x"def80c51",
  2557 => x"0288050d",
  2558 => x"0402f405",
  2559 => x"0d747678",
  2560 => x"53545280",
  2561 => x"71259738",
  2562 => x"72708105",
  2563 => x"5480f52d",
  2564 => x"72708105",
  2565 => x"5481b72d",
  2566 => x"ff115170",
  2567 => x"eb388072",
  2568 => x"81b72d02",
  2569 => x"8c050d04",
  2570 => x"02e8050d",
  2571 => x"77568070",
  2572 => x"56547376",
  2573 => x"24b73880",
  2574 => x"e5f80874",
  2575 => x"2eaf3873",
  2576 => x"5180c9f1",
  2577 => x"2d80def8",
  2578 => x"0880def8",
  2579 => x"08098105",
  2580 => x"7080def8",
  2581 => x"08079f2a",
  2582 => x"77058117",
  2583 => x"57575353",
  2584 => x"74762489",
  2585 => x"3880e5f8",
  2586 => x"087426d3",
  2587 => x"387280de",
  2588 => x"f80c0298",
  2589 => x"050d0402",
  2590 => x"f0050d80",
  2591 => x"def40816",
  2592 => x"5180d0a8",
  2593 => x"2d80def8",
  2594 => x"08802ea0",
  2595 => x"388b5380",
  2596 => x"def80852",
  2597 => x"80e3e851",
  2598 => x"80cff92d",
  2599 => x"80e6a408",
  2600 => x"5473802e",
  2601 => x"873880e3",
  2602 => x"e851732d",
  2603 => x"0290050d",
  2604 => x"0402dc05",
  2605 => x"0d80705a",
  2606 => x"557480de",
  2607 => x"f40825b5",
  2608 => x"3880e5f8",
  2609 => x"08752ead",
  2610 => x"38785180",
  2611 => x"c9f12d80",
  2612 => x"def80809",
  2613 => x"81057080",
  2614 => x"def80807",
  2615 => x"9f2a7605",
  2616 => x"811b5b56",
  2617 => x"547480de",
  2618 => x"f4082589",
  2619 => x"3880e5f8",
  2620 => x"087926d5",
  2621 => x"38805578",
  2622 => x"80e5f808",
  2623 => x"2781e438",
  2624 => x"785180c9",
  2625 => x"f12d80de",
  2626 => x"f808802e",
  2627 => x"81b43880",
  2628 => x"def8088b",
  2629 => x"0580f52d",
  2630 => x"70842a70",
  2631 => x"81067710",
  2632 => x"78842b80",
  2633 => x"e3e80b80",
  2634 => x"f52d5c5c",
  2635 => x"53515556",
  2636 => x"73802e80",
  2637 => x"ce387416",
  2638 => x"822b80d4",
  2639 => x"870b80dd",
  2640 => x"a8120c54",
  2641 => x"77753110",
  2642 => x"80e6a811",
  2643 => x"55569074",
  2644 => x"70810556",
  2645 => x"81b72da0",
  2646 => x"7481b72d",
  2647 => x"7681ff06",
  2648 => x"81165854",
  2649 => x"73802e8b",
  2650 => x"389c5380",
  2651 => x"e3e85280",
  2652 => x"d2fa048b",
  2653 => x"5380def8",
  2654 => x"085280e6",
  2655 => x"aa165180",
  2656 => x"d3b80474",
  2657 => x"16822b80",
  2658 => x"d0f70b80",
  2659 => x"dda8120c",
  2660 => x"547681ff",
  2661 => x"06811658",
  2662 => x"5473802e",
  2663 => x"8b389c53",
  2664 => x"80e3e852",
  2665 => x"80d3af04",
  2666 => x"8b5380de",
  2667 => x"f8085277",
  2668 => x"75311080",
  2669 => x"e6a80551",
  2670 => x"765580cf",
  2671 => x"f92d80d3",
  2672 => x"d7047490",
  2673 => x"29753170",
  2674 => x"1080e6a8",
  2675 => x"05515480",
  2676 => x"def80874",
  2677 => x"81b72d81",
  2678 => x"1959748b",
  2679 => x"24a43880",
  2680 => x"d1f70474",
  2681 => x"90297531",
  2682 => x"701080e6",
  2683 => x"a8058c77",
  2684 => x"31575154",
  2685 => x"807481b7",
  2686 => x"2d9e14ff",
  2687 => x"16565474",
  2688 => x"f33802a4",
  2689 => x"050d0402",
  2690 => x"fc050d80",
  2691 => x"def40813",
  2692 => x"5180d0a8",
  2693 => x"2d80def8",
  2694 => x"08802e8a",
  2695 => x"3880def8",
  2696 => x"085180c1",
  2697 => x"a82d800b",
  2698 => x"80def40c",
  2699 => x"80d1b12d",
  2700 => x"afae2d02",
  2701 => x"84050d04",
  2702 => x"02f4050d",
  2703 => x"7476708c",
  2704 => x"2c708f06",
  2705 => x"80da9408",
  2706 => x"05515353",
  2707 => x"537080f5",
  2708 => x"2d7381b7",
  2709 => x"2d71882c",
  2710 => x"708f0680",
  2711 => x"da940805",
  2712 => x"51517080",
  2713 => x"f52d8114",
  2714 => x"81b72d71",
  2715 => x"842c708f",
  2716 => x"0680da94",
  2717 => x"08055151",
  2718 => x"7080f52d",
  2719 => x"821481b7",
  2720 => x"2d718f06",
  2721 => x"80da9408",
  2722 => x"05527180",
  2723 => x"f52d8314",
  2724 => x"81b72d02",
  2725 => x"8c050d04",
  2726 => x"02f4050d",
  2727 => x"745372fd",
  2728 => x"2eb23872",
  2729 => x"fd248b38",
  2730 => x"72fc2e80",
  2731 => x"d03880d6",
  2732 => x"870472fe",
  2733 => x"2eb93872",
  2734 => x"ff2e0981",
  2735 => x"0680c838",
  2736 => x"80def408",
  2737 => x"5372802e",
  2738 => x"be38ff13",
  2739 => x"80def40c",
  2740 => x"80d68704",
  2741 => x"80def408",
  2742 => x"f4057080",
  2743 => x"def40c53",
  2744 => x"728025a3",
  2745 => x"38800b80",
  2746 => x"def40c80",
  2747 => x"d6870480",
  2748 => x"def40881",
  2749 => x"0580def4",
  2750 => x"0c80d687",
  2751 => x"0480def4",
  2752 => x"088c0580",
  2753 => x"def40c80",
  2754 => x"d1b12d80",
  2755 => x"da805280",
  2756 => x"ded451a2",
  2757 => x"902d80de",
  2758 => x"f4085280",
  2759 => x"ded95180",
  2760 => x"d4b82d80",
  2761 => x"e5f80852",
  2762 => x"80dede51",
  2763 => x"80d4b82d",
  2764 => x"afae2d02",
  2765 => x"8c050d04",
  2766 => x"02fc050d",
  2767 => x"800b80de",
  2768 => x"f40c80d1",
  2769 => x"b12daeaa",
  2770 => x"2d80def8",
  2771 => x"0880dec4",
  2772 => x"0c80dda0",
  2773 => x"51b0d42d",
  2774 => x"0284050d",
  2775 => x"047180e6",
  2776 => x"a40c0400",
  2777 => x"00ffffff",
  2778 => x"ff00ffff",
  2779 => x"ffff00ff",
  2780 => x"ffffff00",
  2781 => x"30313233",
  2782 => x"34353637",
  2783 => x"38394142",
  2784 => x"43444546",
  2785 => x"00000000",
  2786 => x"52657365",
  2787 => x"74000000",
  2788 => x"5363616e",
  2789 => x"6c696e65",
  2790 => x"73000000",
  2791 => x"50414c20",
  2792 => x"2f204e54",
  2793 => x"53430000",
  2794 => x"436f6c6f",
  2795 => x"72000000",
  2796 => x"44696666",
  2797 => x"6963756c",
  2798 => x"74792041",
  2799 => x"00000000",
  2800 => x"44696666",
  2801 => x"6963756c",
  2802 => x"74792042",
  2803 => x"00000000",
  2804 => x"2a537570",
  2805 => x"65726368",
  2806 => x"69702069",
  2807 => x"6e206361",
  2808 => x"72747269",
  2809 => x"64676500",
  2810 => x"2a42616e",
  2811 => x"6b204530",
  2812 => x"00000000",
  2813 => x"2a42616e",
  2814 => x"6b204537",
  2815 => x"00000000",
  2816 => x"53656c65",
  2817 => x"63740000",
  2818 => x"53746172",
  2819 => x"74000000",
  2820 => x"4c6f6164",
  2821 => x"20524f4d",
  2822 => x"20100000",
  2823 => x"45786974",
  2824 => x"00000000",
  2825 => x"524f4d20",
  2826 => x"6c6f6164",
  2827 => x"696e6720",
  2828 => x"6661696c",
  2829 => x"65640000",
  2830 => x"4f4b0000",
  2831 => x"496e6974",
  2832 => x"69616c69",
  2833 => x"7a696e67",
  2834 => x"20534420",
  2835 => x"63617264",
  2836 => x"0a000000",
  2837 => x"16200000",
  2838 => x"14200000",
  2839 => x"15200000",
  2840 => x"53442069",
  2841 => x"6e69742e",
  2842 => x"2e2e0a00",
  2843 => x"53442063",
  2844 => x"61726420",
  2845 => x"72657365",
  2846 => x"74206661",
  2847 => x"696c6564",
  2848 => x"210a0000",
  2849 => x"53444843",
  2850 => x"20657272",
  2851 => x"6f72210a",
  2852 => x"00000000",
  2853 => x"57726974",
  2854 => x"65206661",
  2855 => x"696c6564",
  2856 => x"0a000000",
  2857 => x"52656164",
  2858 => x"20666169",
  2859 => x"6c65640a",
  2860 => x"00000000",
  2861 => x"43617264",
  2862 => x"20696e69",
  2863 => x"74206661",
  2864 => x"696c6564",
  2865 => x"0a000000",
  2866 => x"46415431",
  2867 => x"36202020",
  2868 => x"00000000",
  2869 => x"46415433",
  2870 => x"32202020",
  2871 => x"00000000",
  2872 => x"4e6f2070",
  2873 => x"61727469",
  2874 => x"74696f6e",
  2875 => x"20736967",
  2876 => x"0a000000",
  2877 => x"42616420",
  2878 => x"70617274",
  2879 => x"0a000000",
  2880 => x"4261636b",
  2881 => x"207a7a7a",
  2882 => x"7a207878",
  2883 => x"78780000",
  2884 => x"00000002",
  2885 => x"00002b74",
  2886 => x"00000002",
  2887 => x"00002b88",
  2888 => x"0000035a",
  2889 => x"00000001",
  2890 => x"00002b90",
  2891 => x"00000000",
  2892 => x"00000001",
  2893 => x"00002b9c",
  2894 => x"00000001",
  2895 => x"00000001",
  2896 => x"00002ba8",
  2897 => x"00000002",
  2898 => x"00000001",
  2899 => x"00002bb0",
  2900 => x"00000003",
  2901 => x"00000001",
  2902 => x"00002bc0",
  2903 => x"00000004",
  2904 => x"00000001",
  2905 => x"00002bd0",
  2906 => x"00000005",
  2907 => x"00000001",
  2908 => x"00002be8",
  2909 => x"00000008",
  2910 => x"00000001",
  2911 => x"00002bf4",
  2912 => x"00000009",
  2913 => x"00000002",
  2914 => x"00002c00",
  2915 => x"0000036e",
  2916 => x"00000002",
  2917 => x"00002c08",
  2918 => x"00000a3f",
  2919 => x"00000002",
  2920 => x"00002c10",
  2921 => x"00002b38",
  2922 => x"00000002",
  2923 => x"00002c1c",
  2924 => x"00001747",
  2925 => x"00000000",
  2926 => x"00000000",
  2927 => x"00000000",
  2928 => x"00000004",
  2929 => x"00002c24",
  2930 => x"00002dc0",
  2931 => x"00000004",
  2932 => x"00002c38",
  2933 => x"00002d18",
  2934 => x"00000000",
  2935 => x"00000000",
  2936 => x"00000000",
  2937 => x"00000000",
  2938 => x"00000000",
  2939 => x"00000000",
  2940 => x"00000000",
  2941 => x"00000000",
  2942 => x"00000000",
  2943 => x"00000000",
  2944 => x"00000000",
  2945 => x"00000000",
  2946 => x"00000000",
  2947 => x"00000000",
  2948 => x"00000000",
  2949 => x"00000000",
  2950 => x"00000000",
  2951 => x"00000000",
  2952 => x"00000000",
  2953 => x"761c1c1c",
  2954 => x"1c1c051c",
  2955 => x"1c1c1c1c",
  2956 => x"f2f5fafd",
  2957 => x"5a000000",
  2958 => x"00000000",
  2959 => x"00000000",
  2960 => x"00000000",
  2961 => x"00000000",
  2962 => x"00000000",
  2963 => x"00000000",
  2964 => x"00000000",
  2965 => x"00000000",
  2966 => x"00000000",
  2967 => x"00000000",
  2968 => x"00000000",
  2969 => x"00000000",
  2970 => x"00000000",
  2971 => x"00000000",
  2972 => x"00000000",
  2973 => x"00000000",
  2974 => x"00000000",
  2975 => x"00000000",
  2976 => x"0001ffff",
  2977 => x"0001ffff",
  2978 => x"0001ffff",
  2979 => x"00000000",
  2980 => x"00000000",
  2981 => x"00000004",
  2982 => x"00000000",
  2983 => x"00000000",
  2984 => x"00000002",
  2985 => x"00003328",
  2986 => x"00002877",
  2987 => x"00000002",
  2988 => x"00003346",
  2989 => x"00002877",
  2990 => x"00000002",
  2991 => x"00003364",
  2992 => x"00002877",
  2993 => x"00000002",
  2994 => x"00003382",
  2995 => x"00002877",
  2996 => x"00000002",
  2997 => x"000033a0",
  2998 => x"00002877",
  2999 => x"00000002",
  3000 => x"000033be",
  3001 => x"00002877",
  3002 => x"00000002",
  3003 => x"000033dc",
  3004 => x"00002877",
  3005 => x"00000002",
  3006 => x"000033fa",
  3007 => x"00002877",
  3008 => x"00000002",
  3009 => x"00003418",
  3010 => x"00002877",
  3011 => x"00000002",
  3012 => x"00003436",
  3013 => x"00002877",
  3014 => x"00000002",
  3015 => x"00003454",
  3016 => x"00002877",
  3017 => x"00000002",
  3018 => x"00003472",
  3019 => x"00002877",
  3020 => x"00000002",
  3021 => x"00003490",
  3022 => x"00002877",
  3023 => x"00000004",
  3024 => x"00002f54",
  3025 => x"00000000",
  3026 => x"00000000",
  3027 => x"00000000",
  3028 => x"00002a98",
  3029 => x"4261636b",
  3030 => x"00000000",
  3031 => x"00000000",
  3032 => x"00000000",
  3033 => x"00000000",
  3034 => x"00000000",
  3035 => x"00000000",
  3036 => x"00000000",
  3037 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

