-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80db",
     9 => x"e8080b0b",
    10 => x"80dbec08",
    11 => x"0b0b80db",
    12 => x"f0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"dbf00c0b",
    16 => x"0b80dbec",
    17 => x"0c0b0b80",
    18 => x"dbe80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d4c4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80dbe870",
    57 => x"80e7a827",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a5ed",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80db",
    65 => x"f80c9f0b",
    66 => x"80dbfc0c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"dbfc08ff",
    70 => x"0580dbfc",
    71 => x"0c80dbfc",
    72 => x"088025e8",
    73 => x"3880dbf8",
    74 => x"08ff0580",
    75 => x"dbf80c80",
    76 => x"dbf80880",
    77 => x"25d03880",
    78 => x"0b80dbfc",
    79 => x"0c800b80",
    80 => x"dbf80c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80dbf808",
   100 => x"25913882",
   101 => x"c82d80db",
   102 => x"f808ff05",
   103 => x"80dbf80c",
   104 => x"838a0480",
   105 => x"dbf80880",
   106 => x"dbfc0853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80dbf808",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"dbfc0881",
   116 => x"0580dbfc",
   117 => x"0c80dbfc",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80dbfc",
   121 => x"0c80dbf8",
   122 => x"08810580",
   123 => x"dbf80c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480db",
   128 => x"fc088105",
   129 => x"80dbfc0c",
   130 => x"80dbfc08",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80dbfc",
   134 => x"0c80dbf8",
   135 => x"08810580",
   136 => x"dbf80c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"dc800cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"dc800c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280dc",
   177 => x"80088407",
   178 => x"80dc800c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80d7",
   183 => x"e80c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80dc80",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80db",
   208 => x"e80c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02f8050d",
  1093 => x"028f0580",
  1094 => x"f52d80d7",
  1095 => x"f0085252",
  1096 => x"7080dd95",
  1097 => x"279a3871",
  1098 => x"7181b72d",
  1099 => x"80d7f008",
  1100 => x"810580d7",
  1101 => x"f00c80d7",
  1102 => x"f0085180",
  1103 => x"7181b72d",
  1104 => x"0288050d",
  1105 => x"0402f405",
  1106 => x"0d747084",
  1107 => x"2a708f06",
  1108 => x"80d7ec08",
  1109 => x"057080f5",
  1110 => x"2d545153",
  1111 => x"53a2902d",
  1112 => x"728f0680",
  1113 => x"d7ec0805",
  1114 => x"7080f52d",
  1115 => x"5253a290",
  1116 => x"2d028c05",
  1117 => x"0d0402f4",
  1118 => x"050d7476",
  1119 => x"54527270",
  1120 => x"81055480",
  1121 => x"f52d5170",
  1122 => x"72708105",
  1123 => x"5481b72d",
  1124 => x"70ec3870",
  1125 => x"7281b72d",
  1126 => x"028c050d",
  1127 => x"0402d005",
  1128 => x"0d800b80",
  1129 => x"daa40881",
  1130 => x"8006715d",
  1131 => x"5d59810b",
  1132 => x"ec0c840b",
  1133 => x"ec0c7d52",
  1134 => x"80dc8451",
  1135 => x"80cb912d",
  1136 => x"80dbe808",
  1137 => x"792e80ff",
  1138 => x"3880dc88",
  1139 => x"0879ff12",
  1140 => x"57595774",
  1141 => x"792e8b38",
  1142 => x"81187581",
  1143 => x"2a565874",
  1144 => x"f738f718",
  1145 => x"58815980",
  1146 => x"772580db",
  1147 => x"38775274",
  1148 => x"5184a82d",
  1149 => x"80dde052",
  1150 => x"80dc8451",
  1151 => x"80cde52d",
  1152 => x"80dbe808",
  1153 => x"802ea638",
  1154 => x"80dde05a",
  1155 => x"7ba73883",
  1156 => x"ff567970",
  1157 => x"81055b80",
  1158 => x"f52d7b81",
  1159 => x"1d5de40c",
  1160 => x"e80cff16",
  1161 => x"56758025",
  1162 => x"e938a4b5",
  1163 => x"0480dbe8",
  1164 => x"08598480",
  1165 => x"5780dc84",
  1166 => x"5180cdb4",
  1167 => x"2dfc8017",
  1168 => x"81165657",
  1169 => x"a3e70480",
  1170 => x"dc8808f8",
  1171 => x"0c810be0",
  1172 => x"0c805186",
  1173 => x"da2d86c7",
  1174 => x"2d78802e",
  1175 => x"883880d7",
  1176 => x"f451a4e9",
  1177 => x"0480d99c",
  1178 => x"51afc02d",
  1179 => x"7880dbe8",
  1180 => x"0c02b005",
  1181 => x"0d0402ec",
  1182 => x"050d80dc",
  1183 => x"d40b80d7",
  1184 => x"f00c80dc",
  1185 => x"d4538073",
  1186 => x"81b72d80",
  1187 => x"d9c00851",
  1188 => x"a2c52dba",
  1189 => x"51a2902d",
  1190 => x"ffb408ff",
  1191 => x"b8087098",
  1192 => x"2a535155",
  1193 => x"a2c52d74",
  1194 => x"902a7081",
  1195 => x"ff065254",
  1196 => x"a2c52d74",
  1197 => x"882a7081",
  1198 => x"ff065254",
  1199 => x"a2c52d74",
  1200 => x"81ff0651",
  1201 => x"a2c52d72",
  1202 => x"5280dc90",
  1203 => x"51a2f62d",
  1204 => x"80d7f451",
  1205 => x"afc02d80",
  1206 => x"d9c00884",
  1207 => x"0580d9c0",
  1208 => x"0c029405",
  1209 => x"0d04800b",
  1210 => x"80d9c00c",
  1211 => x"0402ec05",
  1212 => x"0d840bec",
  1213 => x"0cacfd2d",
  1214 => x"a7e32d81",
  1215 => x"f92d8353",
  1216 => x"ace02d81",
  1217 => x"51858d2d",
  1218 => x"ff135372",
  1219 => x"8025f138",
  1220 => x"840bec0c",
  1221 => x"80d68c51",
  1222 => x"86a02d80",
  1223 => x"c1bb2d80",
  1224 => x"dbe80880",
  1225 => x"2e81a538",
  1226 => x"a39d5180",
  1227 => x"d4bb2d80",
  1228 => x"d6a45280",
  1229 => x"dc9051a2",
  1230 => x"f62d80d7",
  1231 => x"f451afc0",
  1232 => x"2dad9f2d",
  1233 => x"a8b42daf",
  1234 => x"d32d80d8",
  1235 => x"880b80f5",
  1236 => x"2d80daa4",
  1237 => x"08708106",
  1238 => x"55565472",
  1239 => x"802e8538",
  1240 => x"73840754",
  1241 => x"74812a70",
  1242 => x"81065153",
  1243 => x"72802e85",
  1244 => x"38738207",
  1245 => x"5474822a",
  1246 => x"70810651",
  1247 => x"5372802e",
  1248 => x"85387381",
  1249 => x"07547483",
  1250 => x"2a708106",
  1251 => x"51537280",
  1252 => x"2e853873",
  1253 => x"88075474",
  1254 => x"842a7081",
  1255 => x"06515372",
  1256 => x"802e8538",
  1257 => x"73900754",
  1258 => x"74852a70",
  1259 => x"81065153",
  1260 => x"72802e85",
  1261 => x"3873a007",
  1262 => x"5473fc0c",
  1263 => x"865380db",
  1264 => x"e8088338",
  1265 => x"845372ec",
  1266 => x"0ca6c404",
  1267 => x"800b80db",
  1268 => x"e80c0294",
  1269 => x"050d0471",
  1270 => x"980c04ff",
  1271 => x"b00880db",
  1272 => x"e80c0481",
  1273 => x"0bffb00c",
  1274 => x"04800bff",
  1275 => x"b00c0402",
  1276 => x"f8050dff",
  1277 => x"b408709f",
  1278 => x"ff065151",
  1279 => x"7080da94",
  1280 => x"082e8c38",
  1281 => x"7080da94",
  1282 => x"0c800b80",
  1283 => x"da900c80",
  1284 => x"da900851",
  1285 => x"81527087",
  1286 => x"e82e8f38",
  1287 => x"7087e824",
  1288 => x"87387111",
  1289 => x"80da900c",
  1290 => x"80527180",
  1291 => x"dbe80c02",
  1292 => x"88050d04",
  1293 => x"02e0050d",
  1294 => x"a9c20480",
  1295 => x"dbe80881",
  1296 => x"f02e0981",
  1297 => x"068a3881",
  1298 => x"0b80da9c",
  1299 => x"0ca9c204",
  1300 => x"80dbe808",
  1301 => x"81e02e09",
  1302 => x"81068a38",
  1303 => x"810b80da",
  1304 => x"a00ca9c2",
  1305 => x"0480dbe8",
  1306 => x"085280da",
  1307 => x"a008802e",
  1308 => x"893880db",
  1309 => x"e8088180",
  1310 => x"05527184",
  1311 => x"2c728f06",
  1312 => x"535380da",
  1313 => x"9c08802e",
  1314 => x"9a387284",
  1315 => x"2980d9c4",
  1316 => x"05721381",
  1317 => x"712b7009",
  1318 => x"73080673",
  1319 => x"0c515353",
  1320 => x"a9b60472",
  1321 => x"842980d9",
  1322 => x"c4057213",
  1323 => x"83712b72",
  1324 => x"0807720c",
  1325 => x"5353800b",
  1326 => x"80daa00c",
  1327 => x"800b80da",
  1328 => x"9c0c80dd",
  1329 => x"9851abd3",
  1330 => x"2d80dbe8",
  1331 => x"08ff24fe",
  1332 => x"ea38a7ef",
  1333 => x"2d80dbe8",
  1334 => x"08802e80",
  1335 => x"ff388156",
  1336 => x"800b80da",
  1337 => x"980880da",
  1338 => x"940880da",
  1339 => x"9c085759",
  1340 => x"59557776",
  1341 => x"06777706",
  1342 => x"54527173",
  1343 => x"2e80c438",
  1344 => x"7280da84",
  1345 => x"1680f52d",
  1346 => x"70842c71",
  1347 => x"8f065255",
  1348 => x"53547380",
  1349 => x"2e9a3872",
  1350 => x"842980d9",
  1351 => x"c4057213",
  1352 => x"81712b70",
  1353 => x"09730806",
  1354 => x"730c5153",
  1355 => x"53aac304",
  1356 => x"72842980",
  1357 => x"d9c40572",
  1358 => x"1383712b",
  1359 => x"72080772",
  1360 => x"0c535375",
  1361 => x"10811656",
  1362 => x"568b7525",
  1363 => x"ffa43873",
  1364 => x"80da9c0c",
  1365 => x"80da9408",
  1366 => x"80da980c",
  1367 => x"800b80db",
  1368 => x"e80c02a0",
  1369 => x"050d0402",
  1370 => x"f8050d80",
  1371 => x"d9c4528f",
  1372 => x"51807270",
  1373 => x"8405540c",
  1374 => x"ff115170",
  1375 => x"8025f238",
  1376 => x"0288050d",
  1377 => x"0402f005",
  1378 => x"0d7551a7",
  1379 => x"e92d7082",
  1380 => x"2cfc0680",
  1381 => x"d9c41172",
  1382 => x"109e0671",
  1383 => x"0870722a",
  1384 => x"70830682",
  1385 => x"742b7009",
  1386 => x"7406760c",
  1387 => x"54515657",
  1388 => x"535153a7",
  1389 => x"e32d7180",
  1390 => x"dbe80c02",
  1391 => x"90050d04",
  1392 => x"02fc050d",
  1393 => x"72518071",
  1394 => x"0c800b84",
  1395 => x"120c0284",
  1396 => x"050d0402",
  1397 => x"f0050d75",
  1398 => x"70088412",
  1399 => x"08535353",
  1400 => x"ff547171",
  1401 => x"2ea838a7",
  1402 => x"e92d8413",
  1403 => x"08708429",
  1404 => x"14881170",
  1405 => x"087081ff",
  1406 => x"06841808",
  1407 => x"81118706",
  1408 => x"841a0c53",
  1409 => x"51555151",
  1410 => x"51a7e32d",
  1411 => x"71547380",
  1412 => x"dbe80c02",
  1413 => x"90050d04",
  1414 => x"02f8050d",
  1415 => x"a7e92de0",
  1416 => x"08708b2a",
  1417 => x"70810651",
  1418 => x"52527080",
  1419 => x"2ea13880",
  1420 => x"dd980870",
  1421 => x"842980dd",
  1422 => x"a0057381",
  1423 => x"ff06710c",
  1424 => x"515180dd",
  1425 => x"98088111",
  1426 => x"870680dd",
  1427 => x"980c5180",
  1428 => x"0b80ddc0",
  1429 => x"0ca7db2d",
  1430 => x"a7e32d02",
  1431 => x"88050d04",
  1432 => x"02fc050d",
  1433 => x"a7e92d81",
  1434 => x"0b80ddc0",
  1435 => x"0ca7e32d",
  1436 => x"80ddc008",
  1437 => x"5170f938",
  1438 => x"0284050d",
  1439 => x"0402fc05",
  1440 => x"0d80dd98",
  1441 => x"51abc02d",
  1442 => x"aae72dac",
  1443 => x"9851a7d7",
  1444 => x"2d028405",
  1445 => x"0d0480dd",
  1446 => x"cc0880db",
  1447 => x"e80c0402",
  1448 => x"fc050d81",
  1449 => x"0b80daa8",
  1450 => x"0c815185",
  1451 => x"8d2d0284",
  1452 => x"050d0402",
  1453 => x"fc050dad",
  1454 => x"bd04a8b4",
  1455 => x"2d80f651",
  1456 => x"ab852d80",
  1457 => x"dbe808f2",
  1458 => x"3880da51",
  1459 => x"ab852d80",
  1460 => x"dbe808e6",
  1461 => x"3880dbe8",
  1462 => x"0880daa8",
  1463 => x"0c80dbe8",
  1464 => x"0851858d",
  1465 => x"2d028405",
  1466 => x"0d0402ec",
  1467 => x"050d7654",
  1468 => x"8052870b",
  1469 => x"881580f5",
  1470 => x"2d565374",
  1471 => x"72248338",
  1472 => x"a0537251",
  1473 => x"83842d81",
  1474 => x"128b1580",
  1475 => x"f52d5452",
  1476 => x"727225de",
  1477 => x"38029405",
  1478 => x"0d0402f0",
  1479 => x"050d80dd",
  1480 => x"cc085481",
  1481 => x"f92d800b",
  1482 => x"80ddd00c",
  1483 => x"7308802e",
  1484 => x"81893882",
  1485 => x"0b80dbfc",
  1486 => x"0c80ddd0",
  1487 => x"088f0680",
  1488 => x"dbf80c73",
  1489 => x"08527183",
  1490 => x"2e963871",
  1491 => x"83268938",
  1492 => x"71812eb0",
  1493 => x"38afa404",
  1494 => x"71852ea0",
  1495 => x"38afa404",
  1496 => x"881480f5",
  1497 => x"2d841508",
  1498 => x"80d6b453",
  1499 => x"545286a0",
  1500 => x"2d718429",
  1501 => x"13700852",
  1502 => x"52afa804",
  1503 => x"7351adea",
  1504 => x"2dafa404",
  1505 => x"80daa408",
  1506 => x"8815082c",
  1507 => x"70810651",
  1508 => x"5271802e",
  1509 => x"883880d6",
  1510 => x"b851afa1",
  1511 => x"0480d6bc",
  1512 => x"5186a02d",
  1513 => x"84140851",
  1514 => x"86a02d80",
  1515 => x"ddd00881",
  1516 => x"0580ddd0",
  1517 => x"0c8c1454",
  1518 => x"aeac0402",
  1519 => x"90050d04",
  1520 => x"7180ddcc",
  1521 => x"0cae9a2d",
  1522 => x"80ddd008",
  1523 => x"ff0580dd",
  1524 => x"d40c0402",
  1525 => x"e8050d80",
  1526 => x"ddcc0880",
  1527 => x"ddd80857",
  1528 => x"5580f651",
  1529 => x"ab852d80",
  1530 => x"dbe80881",
  1531 => x"2a708106",
  1532 => x"51527180",
  1533 => x"2ea438af",
  1534 => x"fd04a8b4",
  1535 => x"2d80f651",
  1536 => x"ab852d80",
  1537 => x"dbe808f2",
  1538 => x"3880daa8",
  1539 => x"08813270",
  1540 => x"80daa80c",
  1541 => x"70525285",
  1542 => x"8d2d800b",
  1543 => x"80ddc40c",
  1544 => x"800b80dd",
  1545 => x"c80c80da",
  1546 => x"a808838d",
  1547 => x"3880da51",
  1548 => x"ab852d80",
  1549 => x"dbe80880",
  1550 => x"2e8c3880",
  1551 => x"ddc40881",
  1552 => x"800780dd",
  1553 => x"c40c80d9",
  1554 => x"51ab852d",
  1555 => x"80dbe808",
  1556 => x"802e8c38",
  1557 => x"80ddc408",
  1558 => x"80c00780",
  1559 => x"ddc40c81",
  1560 => x"9451ab85",
  1561 => x"2d80dbe8",
  1562 => x"08802e8b",
  1563 => x"3880ddc4",
  1564 => x"08900780",
  1565 => x"ddc40c81",
  1566 => x"9151ab85",
  1567 => x"2d80dbe8",
  1568 => x"08802e8b",
  1569 => x"3880ddc4",
  1570 => x"08a00780",
  1571 => x"ddc40c81",
  1572 => x"f551ab85",
  1573 => x"2d80dbe8",
  1574 => x"08802e8b",
  1575 => x"3880ddc4",
  1576 => x"08810780",
  1577 => x"ddc40c81",
  1578 => x"f251ab85",
  1579 => x"2d80dbe8",
  1580 => x"08802e8b",
  1581 => x"3880ddc4",
  1582 => x"08820780",
  1583 => x"ddc40c81",
  1584 => x"eb51ab85",
  1585 => x"2d80dbe8",
  1586 => x"08802e8b",
  1587 => x"3880ddc4",
  1588 => x"08840780",
  1589 => x"ddc40c81",
  1590 => x"f451ab85",
  1591 => x"2d80dbe8",
  1592 => x"08802e8b",
  1593 => x"3880ddc4",
  1594 => x"08880780",
  1595 => x"ddc40c80",
  1596 => x"d851ab85",
  1597 => x"2d80dbe8",
  1598 => x"08802e8c",
  1599 => x"3880ddc8",
  1600 => x"08818007",
  1601 => x"80ddc80c",
  1602 => x"9251ab85",
  1603 => x"2d80dbe8",
  1604 => x"08802e8c",
  1605 => x"3880ddc8",
  1606 => x"0880c007",
  1607 => x"80ddc80c",
  1608 => x"9451ab85",
  1609 => x"2d80dbe8",
  1610 => x"08802e8b",
  1611 => x"3880ddc8",
  1612 => x"08900780",
  1613 => x"ddc80c91",
  1614 => x"51ab852d",
  1615 => x"80dbe808",
  1616 => x"802e8b38",
  1617 => x"80ddc808",
  1618 => x"a00780dd",
  1619 => x"c80c9d51",
  1620 => x"ab852d80",
  1621 => x"dbe80880",
  1622 => x"2e8b3880",
  1623 => x"ddc80881",
  1624 => x"0780ddc8",
  1625 => x"0c9b51ab",
  1626 => x"852d80db",
  1627 => x"e808802e",
  1628 => x"8b3880dd",
  1629 => x"c8088207",
  1630 => x"80ddc80c",
  1631 => x"9c51ab85",
  1632 => x"2d80dbe8",
  1633 => x"08802e8b",
  1634 => x"3880ddc8",
  1635 => x"08840780",
  1636 => x"ddc80ca3",
  1637 => x"51ab852d",
  1638 => x"80dbe808",
  1639 => x"802e8b38",
  1640 => x"80ddc808",
  1641 => x"880780dd",
  1642 => x"c80c81fd",
  1643 => x"51ab852d",
  1644 => x"81fa51ab",
  1645 => x"852db98e",
  1646 => x"0481f551",
  1647 => x"ab852d80",
  1648 => x"dbe80881",
  1649 => x"2a708106",
  1650 => x"51527180",
  1651 => x"2eb33880",
  1652 => x"ddd40852",
  1653 => x"71802e8a",
  1654 => x"38ff1280",
  1655 => x"ddd40cb4",
  1656 => x"810480dd",
  1657 => x"d0081080",
  1658 => x"ddd00805",
  1659 => x"70842916",
  1660 => x"51528812",
  1661 => x"08802e89",
  1662 => x"38ff5188",
  1663 => x"12085271",
  1664 => x"2d81f251",
  1665 => x"ab852d80",
  1666 => x"dbe80881",
  1667 => x"2a708106",
  1668 => x"51527180",
  1669 => x"2eb43880",
  1670 => x"ddd008ff",
  1671 => x"1180ddd4",
  1672 => x"08565353",
  1673 => x"7372258a",
  1674 => x"38811480",
  1675 => x"ddd40cb4",
  1676 => x"ca047210",
  1677 => x"13708429",
  1678 => x"16515288",
  1679 => x"1208802e",
  1680 => x"8938fe51",
  1681 => x"88120852",
  1682 => x"712d81fd",
  1683 => x"51ab852d",
  1684 => x"80dbe808",
  1685 => x"812a7081",
  1686 => x"06515271",
  1687 => x"802eb138",
  1688 => x"80ddd408",
  1689 => x"802e8a38",
  1690 => x"800b80dd",
  1691 => x"d40cb590",
  1692 => x"0480ddd0",
  1693 => x"081080dd",
  1694 => x"d0080570",
  1695 => x"84291651",
  1696 => x"52881208",
  1697 => x"802e8938",
  1698 => x"fd518812",
  1699 => x"0852712d",
  1700 => x"81fa51ab",
  1701 => x"852d80db",
  1702 => x"e808812a",
  1703 => x"70810651",
  1704 => x"5271802e",
  1705 => x"b13880dd",
  1706 => x"d008ff11",
  1707 => x"545280dd",
  1708 => x"d4087325",
  1709 => x"89387280",
  1710 => x"ddd40cb5",
  1711 => x"d6047110",
  1712 => x"12708429",
  1713 => x"16515288",
  1714 => x"1208802e",
  1715 => x"8938fc51",
  1716 => x"88120852",
  1717 => x"712d80dd",
  1718 => x"d4087053",
  1719 => x"5473802e",
  1720 => x"8a388c15",
  1721 => x"ff155555",
  1722 => x"b5dd0482",
  1723 => x"0b80dbfc",
  1724 => x"0c718f06",
  1725 => x"80dbf80c",
  1726 => x"81eb51ab",
  1727 => x"852d80db",
  1728 => x"e808812a",
  1729 => x"70810651",
  1730 => x"5271802e",
  1731 => x"ad387408",
  1732 => x"852e0981",
  1733 => x"06a43888",
  1734 => x"1580f52d",
  1735 => x"ff055271",
  1736 => x"881681b7",
  1737 => x"2d71982b",
  1738 => x"52718025",
  1739 => x"8838800b",
  1740 => x"881681b7",
  1741 => x"2d7451ad",
  1742 => x"ea2d81f4",
  1743 => x"51ab852d",
  1744 => x"80dbe808",
  1745 => x"812a7081",
  1746 => x"06515271",
  1747 => x"802eb338",
  1748 => x"7408852e",
  1749 => x"098106aa",
  1750 => x"38881580",
  1751 => x"f52d8105",
  1752 => x"52718816",
  1753 => x"81b72d71",
  1754 => x"81ff068b",
  1755 => x"1680f52d",
  1756 => x"54527272",
  1757 => x"27873872",
  1758 => x"881681b7",
  1759 => x"2d7451ad",
  1760 => x"ea2d80da",
  1761 => x"51ab852d",
  1762 => x"80dbe808",
  1763 => x"812a7081",
  1764 => x"06515271",
  1765 => x"802e81ad",
  1766 => x"3880ddcc",
  1767 => x"0880ddd4",
  1768 => x"08555373",
  1769 => x"802e8a38",
  1770 => x"8c13ff15",
  1771 => x"5553b7a3",
  1772 => x"04720852",
  1773 => x"71822ea6",
  1774 => x"38718226",
  1775 => x"89387181",
  1776 => x"2eaa38b8",
  1777 => x"c5047183",
  1778 => x"2eb43871",
  1779 => x"842e0981",
  1780 => x"0680f238",
  1781 => x"88130851",
  1782 => x"afc02db8",
  1783 => x"c50480dd",
  1784 => x"d4085188",
  1785 => x"13085271",
  1786 => x"2db8c504",
  1787 => x"810b8814",
  1788 => x"082b80da",
  1789 => x"a4083280",
  1790 => x"daa40cb8",
  1791 => x"99048813",
  1792 => x"80f52d81",
  1793 => x"058b1480",
  1794 => x"f52d5354",
  1795 => x"71742483",
  1796 => x"38805473",
  1797 => x"881481b7",
  1798 => x"2dae9a2d",
  1799 => x"b8c50475",
  1800 => x"08802ea4",
  1801 => x"38750851",
  1802 => x"ab852d80",
  1803 => x"dbe80881",
  1804 => x"06527180",
  1805 => x"2e8c3880",
  1806 => x"ddd40851",
  1807 => x"84160852",
  1808 => x"712d8816",
  1809 => x"5675d838",
  1810 => x"8054800b",
  1811 => x"80dbfc0c",
  1812 => x"738f0680",
  1813 => x"dbf80ca0",
  1814 => x"527380dd",
  1815 => x"d4082e09",
  1816 => x"81069938",
  1817 => x"80ddd008",
  1818 => x"ff057432",
  1819 => x"70098105",
  1820 => x"7072079f",
  1821 => x"2a917131",
  1822 => x"51515353",
  1823 => x"71518384",
  1824 => x"2d811454",
  1825 => x"8e7425c2",
  1826 => x"3880daa8",
  1827 => x"08527180",
  1828 => x"dbe80c02",
  1829 => x"98050d04",
  1830 => x"02f4050d",
  1831 => x"d45281ff",
  1832 => x"720c7108",
  1833 => x"5381ff72",
  1834 => x"0c72882b",
  1835 => x"83fe8006",
  1836 => x"72087081",
  1837 => x"ff065152",
  1838 => x"5381ff72",
  1839 => x"0c727107",
  1840 => x"882b7208",
  1841 => x"7081ff06",
  1842 => x"51525381",
  1843 => x"ff720c72",
  1844 => x"7107882b",
  1845 => x"72087081",
  1846 => x"ff067207",
  1847 => x"80dbe80c",
  1848 => x"5253028c",
  1849 => x"050d0402",
  1850 => x"f4050d74",
  1851 => x"767181ff",
  1852 => x"06d40c53",
  1853 => x"5380dddc",
  1854 => x"08853871",
  1855 => x"892b5271",
  1856 => x"982ad40c",
  1857 => x"71902a70",
  1858 => x"81ff06d4",
  1859 => x"0c517188",
  1860 => x"2a7081ff",
  1861 => x"06d40c51",
  1862 => x"7181ff06",
  1863 => x"d40c7290",
  1864 => x"2a7081ff",
  1865 => x"06d40c51",
  1866 => x"d4087081",
  1867 => x"ff065151",
  1868 => x"82b8bf52",
  1869 => x"7081ff2e",
  1870 => x"09810694",
  1871 => x"3881ff0b",
  1872 => x"d40cd408",
  1873 => x"7081ff06",
  1874 => x"ff145451",
  1875 => x"5171e538",
  1876 => x"7080dbe8",
  1877 => x"0c028c05",
  1878 => x"0d0402fc",
  1879 => x"050d81c7",
  1880 => x"5181ff0b",
  1881 => x"d40cff11",
  1882 => x"51708025",
  1883 => x"f4380284",
  1884 => x"050d0402",
  1885 => x"f4050d81",
  1886 => x"ff0bd40c",
  1887 => x"93538052",
  1888 => x"87fc80c1",
  1889 => x"51b9e72d",
  1890 => x"80dbe808",
  1891 => x"8b3881ff",
  1892 => x"0bd40c81",
  1893 => x"53bba104",
  1894 => x"bada2dff",
  1895 => x"135372de",
  1896 => x"387280db",
  1897 => x"e80c028c",
  1898 => x"050d0402",
  1899 => x"ec050d81",
  1900 => x"0b80dddc",
  1901 => x"0c8454d0",
  1902 => x"08708f2a",
  1903 => x"70810651",
  1904 => x"515372f3",
  1905 => x"3872d00c",
  1906 => x"bada2d80",
  1907 => x"d6c05186",
  1908 => x"a02dd008",
  1909 => x"708f2a70",
  1910 => x"81065151",
  1911 => x"5372f338",
  1912 => x"810bd00c",
  1913 => x"b1538052",
  1914 => x"84d480c0",
  1915 => x"51b9e72d",
  1916 => x"80dbe808",
  1917 => x"812e9338",
  1918 => x"72822ebf",
  1919 => x"38ff1353",
  1920 => x"72e438ff",
  1921 => x"145473ff",
  1922 => x"ae38bada",
  1923 => x"2d83aa52",
  1924 => x"849c80c8",
  1925 => x"51b9e72d",
  1926 => x"80dbe808",
  1927 => x"812e0981",
  1928 => x"069338b9",
  1929 => x"982d80db",
  1930 => x"e80883ff",
  1931 => x"ff065372",
  1932 => x"83aa2e9f",
  1933 => x"38baf32d",
  1934 => x"bcce0480",
  1935 => x"d6cc5186",
  1936 => x"a02d8053",
  1937 => x"bea30480",
  1938 => x"d6e45186",
  1939 => x"a02d8054",
  1940 => x"bdf40481",
  1941 => x"ff0bd40c",
  1942 => x"b154bada",
  1943 => x"2d8fcf53",
  1944 => x"805287fc",
  1945 => x"80f751b9",
  1946 => x"e72d80db",
  1947 => x"e8085580",
  1948 => x"dbe80881",
  1949 => x"2e098106",
  1950 => x"9c3881ff",
  1951 => x"0bd40c82",
  1952 => x"0a52849c",
  1953 => x"80e951b9",
  1954 => x"e72d80db",
  1955 => x"e808802e",
  1956 => x"8d38bada",
  1957 => x"2dff1353",
  1958 => x"72c638bd",
  1959 => x"e70481ff",
  1960 => x"0bd40c80",
  1961 => x"dbe80852",
  1962 => x"87fc80fa",
  1963 => x"51b9e72d",
  1964 => x"80dbe808",
  1965 => x"b23881ff",
  1966 => x"0bd40cd4",
  1967 => x"085381ff",
  1968 => x"0bd40c81",
  1969 => x"ff0bd40c",
  1970 => x"81ff0bd4",
  1971 => x"0c81ff0b",
  1972 => x"d40c7286",
  1973 => x"2a708106",
  1974 => x"76565153",
  1975 => x"72963880",
  1976 => x"dbe80854",
  1977 => x"bdf40473",
  1978 => x"822efedb",
  1979 => x"38ff1454",
  1980 => x"73fee738",
  1981 => x"7380dddc",
  1982 => x"0c738b38",
  1983 => x"815287fc",
  1984 => x"80d051b9",
  1985 => x"e72d81ff",
  1986 => x"0bd40cd0",
  1987 => x"08708f2a",
  1988 => x"70810651",
  1989 => x"515372f3",
  1990 => x"3872d00c",
  1991 => x"81ff0bd4",
  1992 => x"0c815372",
  1993 => x"80dbe80c",
  1994 => x"0294050d",
  1995 => x"0402e805",
  1996 => x"0d785580",
  1997 => x"5681ff0b",
  1998 => x"d40cd008",
  1999 => x"708f2a70",
  2000 => x"81065151",
  2001 => x"5372f338",
  2002 => x"82810bd0",
  2003 => x"0c81ff0b",
  2004 => x"d40c7752",
  2005 => x"87fc80d1",
  2006 => x"51b9e72d",
  2007 => x"80dbc6df",
  2008 => x"5480dbe8",
  2009 => x"08802e8b",
  2010 => x"3880d784",
  2011 => x"5186a02d",
  2012 => x"bfc70481",
  2013 => x"ff0bd40c",
  2014 => x"d4087081",
  2015 => x"ff065153",
  2016 => x"7281fe2e",
  2017 => x"0981069e",
  2018 => x"3880ff53",
  2019 => x"b9982d80",
  2020 => x"dbe80875",
  2021 => x"70840557",
  2022 => x"0cff1353",
  2023 => x"728025ec",
  2024 => x"388156bf",
  2025 => x"ac04ff14",
  2026 => x"5473c838",
  2027 => x"81ff0bd4",
  2028 => x"0c81ff0b",
  2029 => x"d40cd008",
  2030 => x"708f2a70",
  2031 => x"81065151",
  2032 => x"5372f338",
  2033 => x"72d00c75",
  2034 => x"80dbe80c",
  2035 => x"0298050d",
  2036 => x"0402e805",
  2037 => x"0d77797b",
  2038 => x"58555580",
  2039 => x"53727625",
  2040 => x"a4387470",
  2041 => x"81055680",
  2042 => x"f52d7470",
  2043 => x"81055680",
  2044 => x"f52d5252",
  2045 => x"71712e87",
  2046 => x"38815180",
  2047 => x"c0870481",
  2048 => x"1353bfdd",
  2049 => x"04805170",
  2050 => x"80dbe80c",
  2051 => x"0298050d",
  2052 => x"0402ec05",
  2053 => x"0d765574",
  2054 => x"802e80c4",
  2055 => x"389a1580",
  2056 => x"e02d5180",
  2057 => x"cebf2d80",
  2058 => x"dbe80880",
  2059 => x"dbe80880",
  2060 => x"e4900c80",
  2061 => x"dbe80854",
  2062 => x"5480e3ec",
  2063 => x"08802e9b",
  2064 => x"38941580",
  2065 => x"e02d5180",
  2066 => x"cebf2d80",
  2067 => x"dbe80890",
  2068 => x"2b83fff0",
  2069 => x"0a067075",
  2070 => x"07515372",
  2071 => x"80e4900c",
  2072 => x"80e49008",
  2073 => x"5372802e",
  2074 => x"9e3880e3",
  2075 => x"e408fe14",
  2076 => x"712980e3",
  2077 => x"f8080580",
  2078 => x"e4940c70",
  2079 => x"842b80e3",
  2080 => x"f00c5480",
  2081 => x"c1b60480",
  2082 => x"e3fc0880",
  2083 => x"e4900c80",
  2084 => x"e4800880",
  2085 => x"e4940c80",
  2086 => x"e3ec0880",
  2087 => x"2e8c3880",
  2088 => x"e3e40884",
  2089 => x"2b5380c1",
  2090 => x"b10480e4",
  2091 => x"8408842b",
  2092 => x"537280e3",
  2093 => x"f00c0294",
  2094 => x"050d0402",
  2095 => x"d8050d80",
  2096 => x"0b80e3ec",
  2097 => x"0c8454bb",
  2098 => x"ab2d80db",
  2099 => x"e808802e",
  2100 => x"983880dd",
  2101 => x"e0528051",
  2102 => x"bead2d80",
  2103 => x"dbe80880",
  2104 => x"2e8738fe",
  2105 => x"5480c1f1",
  2106 => x"04ff1454",
  2107 => x"738024d7",
  2108 => x"38738e38",
  2109 => x"80d79451",
  2110 => x"86a02d73",
  2111 => x"5580c7cf",
  2112 => x"04805681",
  2113 => x"0b80e498",
  2114 => x"0c885380",
  2115 => x"d7a85280",
  2116 => x"de9651bf",
  2117 => x"d12d80db",
  2118 => x"e808762e",
  2119 => x"09810689",
  2120 => x"3880dbe8",
  2121 => x"0880e498",
  2122 => x"0c885380",
  2123 => x"d7b45280",
  2124 => x"deb251bf",
  2125 => x"d12d80db",
  2126 => x"e8088938",
  2127 => x"80dbe808",
  2128 => x"80e4980c",
  2129 => x"80e49808",
  2130 => x"802e8184",
  2131 => x"3880e1a6",
  2132 => x"0b80f52d",
  2133 => x"80e1a70b",
  2134 => x"80f52d71",
  2135 => x"982b7190",
  2136 => x"2b0780e1",
  2137 => x"a80b80f5",
  2138 => x"2d70882b",
  2139 => x"720780e1",
  2140 => x"a90b80f5",
  2141 => x"2d710780",
  2142 => x"e1de0b80",
  2143 => x"f52d80e1",
  2144 => x"df0b80f5",
  2145 => x"2d71882b",
  2146 => x"07535f54",
  2147 => x"525a5657",
  2148 => x"557381ab",
  2149 => x"aa2e0981",
  2150 => x"06903875",
  2151 => x"5180ce8e",
  2152 => x"2d80dbe8",
  2153 => x"085680c3",
  2154 => x"b9047382",
  2155 => x"d4d52e89",
  2156 => x"3880d7c0",
  2157 => x"5180c486",
  2158 => x"0480dde0",
  2159 => x"527551be",
  2160 => x"ad2d80db",
  2161 => x"e8085580",
  2162 => x"dbe80880",
  2163 => x"2e848038",
  2164 => x"885380d7",
  2165 => x"b45280de",
  2166 => x"b251bfd1",
  2167 => x"2d80dbe8",
  2168 => x"088b3881",
  2169 => x"0b80e3ec",
  2170 => x"0c80c48d",
  2171 => x"04885380",
  2172 => x"d7a85280",
  2173 => x"de9651bf",
  2174 => x"d12d80db",
  2175 => x"e808802e",
  2176 => x"8c3880d7",
  2177 => x"d45186a0",
  2178 => x"2d80c4ec",
  2179 => x"0480e1de",
  2180 => x"0b80f52d",
  2181 => x"547380d5",
  2182 => x"2e098106",
  2183 => x"80ce3880",
  2184 => x"e1df0b80",
  2185 => x"f52d5473",
  2186 => x"81aa2e09",
  2187 => x"8106bd38",
  2188 => x"800b80dd",
  2189 => x"e00b80f5",
  2190 => x"2d565474",
  2191 => x"81e92e83",
  2192 => x"38815474",
  2193 => x"81eb2e8c",
  2194 => x"38805573",
  2195 => x"752e0981",
  2196 => x"0682fc38",
  2197 => x"80ddeb0b",
  2198 => x"80f52d55",
  2199 => x"748e3880",
  2200 => x"ddec0b80",
  2201 => x"f52d5473",
  2202 => x"822e8738",
  2203 => x"805580c7",
  2204 => x"cf0480dd",
  2205 => x"ed0b80f5",
  2206 => x"2d7080e3",
  2207 => x"e40cff05",
  2208 => x"80e3e80c",
  2209 => x"80ddee0b",
  2210 => x"80f52d80",
  2211 => x"ddef0b80",
  2212 => x"f52d5876",
  2213 => x"05778280",
  2214 => x"29057080",
  2215 => x"e3f40c80",
  2216 => x"ddf00b80",
  2217 => x"f52d7080",
  2218 => x"e4880c80",
  2219 => x"e3ec0859",
  2220 => x"57587680",
  2221 => x"2e81b838",
  2222 => x"885380d7",
  2223 => x"b45280de",
  2224 => x"b251bfd1",
  2225 => x"2d80dbe8",
  2226 => x"08828438",
  2227 => x"80e3e408",
  2228 => x"70842b80",
  2229 => x"e3f00c70",
  2230 => x"80e4840c",
  2231 => x"80de850b",
  2232 => x"80f52d80",
  2233 => x"de840b80",
  2234 => x"f52d7182",
  2235 => x"80290580",
  2236 => x"de860b80",
  2237 => x"f52d7084",
  2238 => x"80802912",
  2239 => x"80de870b",
  2240 => x"80f52d70",
  2241 => x"81800a29",
  2242 => x"127080e4",
  2243 => x"8c0c80e4",
  2244 => x"88087129",
  2245 => x"80e3f408",
  2246 => x"057080e3",
  2247 => x"f80c80de",
  2248 => x"8d0b80f5",
  2249 => x"2d80de8c",
  2250 => x"0b80f52d",
  2251 => x"71828029",
  2252 => x"0580de8e",
  2253 => x"0b80f52d",
  2254 => x"70848080",
  2255 => x"291280de",
  2256 => x"8f0b80f5",
  2257 => x"2d70982b",
  2258 => x"81f00a06",
  2259 => x"72057080",
  2260 => x"e3fc0cfe",
  2261 => x"117e2977",
  2262 => x"0580e480",
  2263 => x"0c525952",
  2264 => x"43545e51",
  2265 => x"5259525d",
  2266 => x"57595780",
  2267 => x"c7c70480",
  2268 => x"ddf20b80",
  2269 => x"f52d80dd",
  2270 => x"f10b80f5",
  2271 => x"2d718280",
  2272 => x"29057080",
  2273 => x"e3f00c70",
  2274 => x"a02983ff",
  2275 => x"0570892a",
  2276 => x"7080e484",
  2277 => x"0c80ddf7",
  2278 => x"0b80f52d",
  2279 => x"80ddf60b",
  2280 => x"80f52d71",
  2281 => x"82802905",
  2282 => x"7080e48c",
  2283 => x"0c7b7129",
  2284 => x"1e7080e4",
  2285 => x"800c7d80",
  2286 => x"e3fc0c73",
  2287 => x"0580e3f8",
  2288 => x"0c555e51",
  2289 => x"51555580",
  2290 => x"5180c091",
  2291 => x"2d815574",
  2292 => x"80dbe80c",
  2293 => x"02a8050d",
  2294 => x"0402ec05",
  2295 => x"0d767087",
  2296 => x"2c7180ff",
  2297 => x"06555654",
  2298 => x"80e3ec08",
  2299 => x"8a387388",
  2300 => x"2c7481ff",
  2301 => x"06545580",
  2302 => x"dde05280",
  2303 => x"e3f40815",
  2304 => x"51bead2d",
  2305 => x"80dbe808",
  2306 => x"5480dbe8",
  2307 => x"08802ebb",
  2308 => x"3880e3ec",
  2309 => x"08802e9c",
  2310 => x"38728429",
  2311 => x"80dde005",
  2312 => x"70085253",
  2313 => x"80ce8e2d",
  2314 => x"80dbe808",
  2315 => x"f00a0653",
  2316 => x"80c8c904",
  2317 => x"721080dd",
  2318 => x"e0057080",
  2319 => x"e02d5253",
  2320 => x"80cebf2d",
  2321 => x"80dbe808",
  2322 => x"53725473",
  2323 => x"80dbe80c",
  2324 => x"0294050d",
  2325 => x"0402e005",
  2326 => x"0d797084",
  2327 => x"2c80e494",
  2328 => x"0805718f",
  2329 => x"06525553",
  2330 => x"728a3880",
  2331 => x"dde05273",
  2332 => x"51bead2d",
  2333 => x"72a02980",
  2334 => x"dde00554",
  2335 => x"807480f5",
  2336 => x"2d565374",
  2337 => x"732e8338",
  2338 => x"81537481",
  2339 => x"e52e81f5",
  2340 => x"38817074",
  2341 => x"06545872",
  2342 => x"802e81e9",
  2343 => x"388b1480",
  2344 => x"f52d7083",
  2345 => x"2a790658",
  2346 => x"56769c38",
  2347 => x"80daac08",
  2348 => x"53728938",
  2349 => x"7280e1e0",
  2350 => x"0b81b72d",
  2351 => x"7680daac",
  2352 => x"0c735380",
  2353 => x"cb870475",
  2354 => x"8f2e0981",
  2355 => x"0681b638",
  2356 => x"749f068d",
  2357 => x"2980e1d3",
  2358 => x"11515381",
  2359 => x"1480f52d",
  2360 => x"73708105",
  2361 => x"5581b72d",
  2362 => x"831480f5",
  2363 => x"2d737081",
  2364 => x"055581b7",
  2365 => x"2d851480",
  2366 => x"f52d7370",
  2367 => x"81055581",
  2368 => x"b72d8714",
  2369 => x"80f52d73",
  2370 => x"70810555",
  2371 => x"81b72d89",
  2372 => x"1480f52d",
  2373 => x"73708105",
  2374 => x"5581b72d",
  2375 => x"8e1480f5",
  2376 => x"2d737081",
  2377 => x"055581b7",
  2378 => x"2d901480",
  2379 => x"f52d7370",
  2380 => x"81055581",
  2381 => x"b72d9214",
  2382 => x"80f52d73",
  2383 => x"70810555",
  2384 => x"81b72d94",
  2385 => x"1480f52d",
  2386 => x"73708105",
  2387 => x"5581b72d",
  2388 => x"961480f5",
  2389 => x"2d737081",
  2390 => x"055581b7",
  2391 => x"2d981480",
  2392 => x"f52d7370",
  2393 => x"81055581",
  2394 => x"b72d9c14",
  2395 => x"80f52d73",
  2396 => x"70810555",
  2397 => x"81b72d9e",
  2398 => x"1480f52d",
  2399 => x"7381b72d",
  2400 => x"7780daac",
  2401 => x"0c805372",
  2402 => x"80dbe80c",
  2403 => x"02a0050d",
  2404 => x"0402cc05",
  2405 => x"0d7e605e",
  2406 => x"5a800b80",
  2407 => x"e4900880",
  2408 => x"e4940859",
  2409 => x"5c568058",
  2410 => x"80e3f008",
  2411 => x"782e81bc",
  2412 => x"38778f06",
  2413 => x"a0175754",
  2414 => x"73913880",
  2415 => x"dde05276",
  2416 => x"51811757",
  2417 => x"bead2d80",
  2418 => x"dde05680",
  2419 => x"7680f52d",
  2420 => x"56547474",
  2421 => x"2e833881",
  2422 => x"547481e5",
  2423 => x"2e818138",
  2424 => x"81707506",
  2425 => x"555c7380",
  2426 => x"2e80f538",
  2427 => x"8b1680f5",
  2428 => x"2d980659",
  2429 => x"7880e938",
  2430 => x"8b537c52",
  2431 => x"7551bfd1",
  2432 => x"2d80dbe8",
  2433 => x"0880d938",
  2434 => x"9c160851",
  2435 => x"80ce8e2d",
  2436 => x"80dbe808",
  2437 => x"841b0c9a",
  2438 => x"1680e02d",
  2439 => x"5180cebf",
  2440 => x"2d80dbe8",
  2441 => x"0880dbe8",
  2442 => x"08881c0c",
  2443 => x"80dbe808",
  2444 => x"555580e3",
  2445 => x"ec08802e",
  2446 => x"9a389416",
  2447 => x"80e02d51",
  2448 => x"80cebf2d",
  2449 => x"80dbe808",
  2450 => x"902b83ff",
  2451 => x"f00a0670",
  2452 => x"16515473",
  2453 => x"881b0c78",
  2454 => x"7a0c7b54",
  2455 => x"80cdaa04",
  2456 => x"81185880",
  2457 => x"e3f00878",
  2458 => x"26fec638",
  2459 => x"80e3ec08",
  2460 => x"802eb538",
  2461 => x"7a5180c7",
  2462 => x"d92d80db",
  2463 => x"e80880db",
  2464 => x"e80880ff",
  2465 => x"fffff806",
  2466 => x"555b7380",
  2467 => x"fffffff8",
  2468 => x"2e963880",
  2469 => x"dbe808fe",
  2470 => x"0580e3e4",
  2471 => x"082980e3",
  2472 => x"f8080557",
  2473 => x"80cba604",
  2474 => x"80547380",
  2475 => x"dbe80c02",
  2476 => x"b4050d04",
  2477 => x"02f4050d",
  2478 => x"74700881",
  2479 => x"05710c70",
  2480 => x"0880e3e8",
  2481 => x"08065353",
  2482 => x"71903888",
  2483 => x"13085180",
  2484 => x"c7d92d80",
  2485 => x"dbe80888",
  2486 => x"140c810b",
  2487 => x"80dbe80c",
  2488 => x"028c050d",
  2489 => x"0402f005",
  2490 => x"0d758811",
  2491 => x"08fe0580",
  2492 => x"e3e40829",
  2493 => x"80e3f808",
  2494 => x"11720880",
  2495 => x"e3e80806",
  2496 => x"05795553",
  2497 => x"5454bead",
  2498 => x"2d029005",
  2499 => x"0d0402f4",
  2500 => x"050d7470",
  2501 => x"882a83fe",
  2502 => x"80067072",
  2503 => x"982a0772",
  2504 => x"882b87fc",
  2505 => x"80800673",
  2506 => x"982b81f0",
  2507 => x"0a067173",
  2508 => x"070780db",
  2509 => x"e80c5651",
  2510 => x"5351028c",
  2511 => x"050d0402",
  2512 => x"f8050d02",
  2513 => x"8e0580f5",
  2514 => x"2d74882b",
  2515 => x"077083ff",
  2516 => x"ff0680db",
  2517 => x"e80c5102",
  2518 => x"88050d04",
  2519 => x"02f4050d",
  2520 => x"74767853",
  2521 => x"54528071",
  2522 => x"25973872",
  2523 => x"70810554",
  2524 => x"80f52d72",
  2525 => x"70810554",
  2526 => x"81b72dff",
  2527 => x"115170eb",
  2528 => x"38807281",
  2529 => x"b72d028c",
  2530 => x"050d0402",
  2531 => x"e8050d77",
  2532 => x"56807056",
  2533 => x"54737624",
  2534 => x"b73880e3",
  2535 => x"f008742e",
  2536 => x"af387351",
  2537 => x"80c8d52d",
  2538 => x"80dbe808",
  2539 => x"80dbe808",
  2540 => x"09810570",
  2541 => x"80dbe808",
  2542 => x"079f2a77",
  2543 => x"05811757",
  2544 => x"57535374",
  2545 => x"76248938",
  2546 => x"80e3f008",
  2547 => x"7426d338",
  2548 => x"7280dbe8",
  2549 => x"0c029805",
  2550 => x"0d0402f0",
  2551 => x"050d80db",
  2552 => x"e4081651",
  2553 => x"80cf8b2d",
  2554 => x"80dbe808",
  2555 => x"802ea038",
  2556 => x"8b5380db",
  2557 => x"e8085280",
  2558 => x"e1e05180",
  2559 => x"cedc2d80",
  2560 => x"e49c0854",
  2561 => x"73802e87",
  2562 => x"3880e1e0",
  2563 => x"51732d02",
  2564 => x"90050d04",
  2565 => x"02dc050d",
  2566 => x"80705a55",
  2567 => x"7480dbe4",
  2568 => x"0825b538",
  2569 => x"80e3f008",
  2570 => x"752ead38",
  2571 => x"785180c8",
  2572 => x"d52d80db",
  2573 => x"e8080981",
  2574 => x"057080db",
  2575 => x"e808079f",
  2576 => x"2a760581",
  2577 => x"1b5b5654",
  2578 => x"7480dbe4",
  2579 => x"08258938",
  2580 => x"80e3f008",
  2581 => x"7926d538",
  2582 => x"80557880",
  2583 => x"e3f00827",
  2584 => x"81e43878",
  2585 => x"5180c8d5",
  2586 => x"2d80dbe8",
  2587 => x"08802e81",
  2588 => x"b43880db",
  2589 => x"e8088b05",
  2590 => x"80f52d70",
  2591 => x"842a7081",
  2592 => x"06771078",
  2593 => x"842b80e1",
  2594 => x"e00b80f5",
  2595 => x"2d5c5c53",
  2596 => x"51555673",
  2597 => x"802e80ce",
  2598 => x"38741682",
  2599 => x"2b80d2ea",
  2600 => x"0b80dab8",
  2601 => x"120c5477",
  2602 => x"75311080",
  2603 => x"e4a01155",
  2604 => x"56907470",
  2605 => x"81055681",
  2606 => x"b72da074",
  2607 => x"81b72d76",
  2608 => x"81ff0681",
  2609 => x"16585473",
  2610 => x"802e8b38",
  2611 => x"9c5380e1",
  2612 => x"e05280d1",
  2613 => x"dd048b53",
  2614 => x"80dbe808",
  2615 => x"5280e4a2",
  2616 => x"165180d2",
  2617 => x"9b047416",
  2618 => x"822b80cf",
  2619 => x"da0b80da",
  2620 => x"b8120c54",
  2621 => x"7681ff06",
  2622 => x"81165854",
  2623 => x"73802e8b",
  2624 => x"389c5380",
  2625 => x"e1e05280",
  2626 => x"d292048b",
  2627 => x"5380dbe8",
  2628 => x"08527775",
  2629 => x"311080e4",
  2630 => x"a0055176",
  2631 => x"5580cedc",
  2632 => x"2d80d2ba",
  2633 => x"04749029",
  2634 => x"75317010",
  2635 => x"80e4a005",
  2636 => x"515480db",
  2637 => x"e8087481",
  2638 => x"b72d8119",
  2639 => x"59748b24",
  2640 => x"a43880d0",
  2641 => x"da047490",
  2642 => x"29753170",
  2643 => x"1080e4a0",
  2644 => x"058c7731",
  2645 => x"57515480",
  2646 => x"7481b72d",
  2647 => x"9e14ff16",
  2648 => x"565474f3",
  2649 => x"3802a405",
  2650 => x"0d0402fc",
  2651 => x"050d80db",
  2652 => x"e4081351",
  2653 => x"80cf8b2d",
  2654 => x"80dbe808",
  2655 => x"802e8a38",
  2656 => x"80dbe808",
  2657 => x"5180c091",
  2658 => x"2d800b80",
  2659 => x"dbe40c80",
  2660 => x"d0942dae",
  2661 => x"9a2d0284",
  2662 => x"050d0402",
  2663 => x"fc050d72",
  2664 => x"5170fd2e",
  2665 => x"b23870fd",
  2666 => x"248b3870",
  2667 => x"fc2e80d0",
  2668 => x"3880d48a",
  2669 => x"0470fe2e",
  2670 => x"b93870ff",
  2671 => x"2e098106",
  2672 => x"80c83880",
  2673 => x"dbe40851",
  2674 => x"70802ebe",
  2675 => x"38ff1180",
  2676 => x"dbe40c80",
  2677 => x"d48a0480",
  2678 => x"dbe408f0",
  2679 => x"057080db",
  2680 => x"e40c5170",
  2681 => x"8025a338",
  2682 => x"800b80db",
  2683 => x"e40c80d4",
  2684 => x"8a0480db",
  2685 => x"e4088105",
  2686 => x"80dbe40c",
  2687 => x"80d48a04",
  2688 => x"80dbe408",
  2689 => x"900580db",
  2690 => x"e40c80d0",
  2691 => x"942dae9a",
  2692 => x"2d028405",
  2693 => x"0d0402fc",
  2694 => x"050d800b",
  2695 => x"80dbe40c",
  2696 => x"80d0942d",
  2697 => x"ad962d80",
  2698 => x"dbe80880",
  2699 => x"dbd40c80",
  2700 => x"dab051af",
  2701 => x"c02d0284",
  2702 => x"050d0471",
  2703 => x"80e49c0c",
  2704 => x"04000000",
  2705 => x"00ffffff",
  2706 => x"ff00ffff",
  2707 => x"ffff00ff",
  2708 => x"ffffff00",
  2709 => x"30313233",
  2710 => x"34353637",
  2711 => x"38394142",
  2712 => x"43444546",
  2713 => x"00000000",
  2714 => x"44656275",
  2715 => x"67000000",
  2716 => x"52657365",
  2717 => x"74000000",
  2718 => x"5363616e",
  2719 => x"6c696e65",
  2720 => x"73000000",
  2721 => x"50414c20",
  2722 => x"2f204e54",
  2723 => x"53430000",
  2724 => x"436f6c6f",
  2725 => x"72000000",
  2726 => x"44696666",
  2727 => x"6963756c",
  2728 => x"74792041",
  2729 => x"00000000",
  2730 => x"44696666",
  2731 => x"6963756c",
  2732 => x"74792042",
  2733 => x"00000000",
  2734 => x"53757065",
  2735 => x"72636869",
  2736 => x"7020696e",
  2737 => x"20636172",
  2738 => x"74726964",
  2739 => x"67650000",
  2740 => x"53656c65",
  2741 => x"63740000",
  2742 => x"53746172",
  2743 => x"74000000",
  2744 => x"4c6f6164",
  2745 => x"20524f4d",
  2746 => x"20100000",
  2747 => x"45786974",
  2748 => x"00000000",
  2749 => x"524f4d20",
  2750 => x"6c6f6164",
  2751 => x"696e6720",
  2752 => x"6661696c",
  2753 => x"65640000",
  2754 => x"4f4b0000",
  2755 => x"496e6974",
  2756 => x"69616c69",
  2757 => x"7a696e67",
  2758 => x"20534420",
  2759 => x"63617264",
  2760 => x"0a000000",
  2761 => x"436f6c6c",
  2762 => x"6563746f",
  2763 => x"72566973",
  2764 => x"696f6e00",
  2765 => x"16200000",
  2766 => x"14200000",
  2767 => x"15200000",
  2768 => x"53442069",
  2769 => x"6e69742e",
  2770 => x"2e2e0a00",
  2771 => x"53442063",
  2772 => x"61726420",
  2773 => x"72657365",
  2774 => x"74206661",
  2775 => x"696c6564",
  2776 => x"210a0000",
  2777 => x"53444843",
  2778 => x"20657272",
  2779 => x"6f72210a",
  2780 => x"00000000",
  2781 => x"57726974",
  2782 => x"65206661",
  2783 => x"696c6564",
  2784 => x"0a000000",
  2785 => x"52656164",
  2786 => x"20666169",
  2787 => x"6c65640a",
  2788 => x"00000000",
  2789 => x"43617264",
  2790 => x"20696e69",
  2791 => x"74206661",
  2792 => x"696c6564",
  2793 => x"0a000000",
  2794 => x"46415431",
  2795 => x"36202020",
  2796 => x"00000000",
  2797 => x"46415433",
  2798 => x"32202020",
  2799 => x"00000000",
  2800 => x"4e6f2070",
  2801 => x"61727469",
  2802 => x"74696f6e",
  2803 => x"20736967",
  2804 => x"0a000000",
  2805 => x"42616420",
  2806 => x"70617274",
  2807 => x"0a000000",
  2808 => x"4261636b",
  2809 => x"00000000",
  2810 => x"00000002",
  2811 => x"00002a54",
  2812 => x"00002e54",
  2813 => x"00000002",
  2814 => x"00002e10",
  2815 => x"000012e6",
  2816 => x"00000002",
  2817 => x"00002a68",
  2818 => x"00001276",
  2819 => x"00000002",
  2820 => x"00002a70",
  2821 => x"0000035a",
  2822 => x"00000001",
  2823 => x"00002a78",
  2824 => x"00000000",
  2825 => x"00000001",
  2826 => x"00002a84",
  2827 => x"00000001",
  2828 => x"00000001",
  2829 => x"00002a90",
  2830 => x"00000002",
  2831 => x"00000001",
  2832 => x"00002a98",
  2833 => x"00000003",
  2834 => x"00000001",
  2835 => x"00002aa8",
  2836 => x"00000004",
  2837 => x"00000001",
  2838 => x"00002ab8",
  2839 => x"00000005",
  2840 => x"00000002",
  2841 => x"00002ad0",
  2842 => x"0000036e",
  2843 => x"00000002",
  2844 => x"00002ad8",
  2845 => x"00000a3f",
  2846 => x"00000002",
  2847 => x"00002ae0",
  2848 => x"00002a16",
  2849 => x"00000002",
  2850 => x"00002aec",
  2851 => x"000016b3",
  2852 => x"00000000",
  2853 => x"00000000",
  2854 => x"00000000",
  2855 => x"00000004",
  2856 => x"00002af4",
  2857 => x"00002c9c",
  2858 => x"00000004",
  2859 => x"00002b08",
  2860 => x"00002bf4",
  2861 => x"00000000",
  2862 => x"00000000",
  2863 => x"00000000",
  2864 => x"00000000",
  2865 => x"00000000",
  2866 => x"00000000",
  2867 => x"00000000",
  2868 => x"00000000",
  2869 => x"00000000",
  2870 => x"00000000",
  2871 => x"00000000",
  2872 => x"00000000",
  2873 => x"00000000",
  2874 => x"00000000",
  2875 => x"00000000",
  2876 => x"00000000",
  2877 => x"00000000",
  2878 => x"00000000",
  2879 => x"00000000",
  2880 => x"00000000",
  2881 => x"76f55a1c",
  2882 => x"f21c1c1c",
  2883 => x"1c1c1c1c",
  2884 => x"00000000",
  2885 => x"00000fff",
  2886 => x"00000fff",
  2887 => x"00000000",
  2888 => x"00000000",
  2889 => x"00000006",
  2890 => x"00000000",
  2891 => x"00000000",
  2892 => x"00000002",
  2893 => x"00003220",
  2894 => x"000027da",
  2895 => x"00000002",
  2896 => x"0000323e",
  2897 => x"000027da",
  2898 => x"00000002",
  2899 => x"0000325c",
  2900 => x"000027da",
  2901 => x"00000002",
  2902 => x"0000327a",
  2903 => x"000027da",
  2904 => x"00000002",
  2905 => x"00003298",
  2906 => x"000027da",
  2907 => x"00000002",
  2908 => x"000032b6",
  2909 => x"000027da",
  2910 => x"00000002",
  2911 => x"000032d4",
  2912 => x"000027da",
  2913 => x"00000002",
  2914 => x"000032f2",
  2915 => x"000027da",
  2916 => x"00000002",
  2917 => x"00003310",
  2918 => x"000027da",
  2919 => x"00000002",
  2920 => x"0000332e",
  2921 => x"000027da",
  2922 => x"00000002",
  2923 => x"0000334c",
  2924 => x"000027da",
  2925 => x"00000002",
  2926 => x"0000336a",
  2927 => x"000027da",
  2928 => x"00000002",
  2929 => x"00003388",
  2930 => x"000027da",
  2931 => x"00000004",
  2932 => x"00002be0",
  2933 => x"00000000",
  2934 => x"00000000",
  2935 => x"00000000",
  2936 => x"0000299b",
  2937 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

