-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80dd",
     9 => x"a0080b0b",
    10 => x"80dda408",
    11 => x"0b0b80dd",
    12 => x"a8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"dda80c0b",
    16 => x"0b80dda4",
    17 => x"0c0b0b80",
    18 => x"dda00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d5b8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80dda070",
    57 => x"80e7d827",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a6b2",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80dd",
    65 => x"b00c9f0b",
    66 => x"80ddb40c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"ddb408ff",
    70 => x"0580ddb4",
    71 => x"0c80ddb4",
    72 => x"088025e8",
    73 => x"3880ddb0",
    74 => x"08ff0580",
    75 => x"ddb00c80",
    76 => x"ddb00880",
    77 => x"25d03880",
    78 => x"0b80ddb4",
    79 => x"0c800b80",
    80 => x"ddb00c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80ddb008",
   100 => x"25913882",
   101 => x"c82d80dd",
   102 => x"b008ff05",
   103 => x"80ddb00c",
   104 => x"838a0480",
   105 => x"ddb00880",
   106 => x"ddb40853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80ddb008",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"ddb40881",
   116 => x"0580ddb4",
   117 => x"0c80ddb4",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80ddb4",
   121 => x"0c80ddb0",
   122 => x"08810580",
   123 => x"ddb00c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480dd",
   128 => x"b4088105",
   129 => x"80ddb40c",
   130 => x"80ddb408",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80ddb4",
   134 => x"0c80ddb0",
   135 => x"08810580",
   136 => x"ddb00c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"ddb80cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"ddb80c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280dd",
   177 => x"b8088407",
   178 => x"80ddb80c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80d8",
   183 => x"dc0c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80ddb8",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80dd",
   208 => x"a00c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02f4050d",
  1093 => x"80d8f40b",
  1094 => x"80f52d80",
  1095 => x"dbdc0870",
  1096 => x"81065354",
  1097 => x"5270802e",
  1098 => x"85387184",
  1099 => x"07527281",
  1100 => x"2a708106",
  1101 => x"51517080",
  1102 => x"2e853871",
  1103 => x"82075272",
  1104 => x"822a7081",
  1105 => x"06515170",
  1106 => x"802e8538",
  1107 => x"71810752",
  1108 => x"72832a70",
  1109 => x"81065151",
  1110 => x"70802e85",
  1111 => x"38718807",
  1112 => x"5272842a",
  1113 => x"70810651",
  1114 => x"5170802e",
  1115 => x"85387190",
  1116 => x"07527285",
  1117 => x"2a708106",
  1118 => x"51517080",
  1119 => x"2e853871",
  1120 => x"a0075272",
  1121 => x"882a7081",
  1122 => x"06515170",
  1123 => x"802e8638",
  1124 => x"7180c007",
  1125 => x"5272892a",
  1126 => x"70810651",
  1127 => x"5170802e",
  1128 => x"86387181",
  1129 => x"80075271",
  1130 => x"fc0c7180",
  1131 => x"dda00c02",
  1132 => x"8c050d04",
  1133 => x"02cc050d",
  1134 => x"7e5d800b",
  1135 => x"80dbdc08",
  1136 => x"81800671",
  1137 => x"5c5d5b81",
  1138 => x"0bec0c84",
  1139 => x"0bec0c7c",
  1140 => x"5280ddbc",
  1141 => x"5180cc86",
  1142 => x"2d80dda0",
  1143 => x"087b2e80",
  1144 => x"ff3880dd",
  1145 => x"c0087bff",
  1146 => x"12575957",
  1147 => x"747b2e8b",
  1148 => x"38811875",
  1149 => x"812a5658",
  1150 => x"74f738f7",
  1151 => x"1858815b",
  1152 => x"80772580",
  1153 => x"db387752",
  1154 => x"745184a8",
  1155 => x"2d80de90",
  1156 => x"5280ddbc",
  1157 => x"5180cedb",
  1158 => x"2d80dda0",
  1159 => x"08802ea6",
  1160 => x"3880de90",
  1161 => x"597ba738",
  1162 => x"83ff5678",
  1163 => x"7081055a",
  1164 => x"80f52d7a",
  1165 => x"811c5ce4",
  1166 => x"0ce80cff",
  1167 => x"16567580",
  1168 => x"25e938a4",
  1169 => x"ce0480dd",
  1170 => x"a0085b84",
  1171 => x"805780dd",
  1172 => x"bc5180ce",
  1173 => x"aa2dfc80",
  1174 => x"17811656",
  1175 => x"57a48004",
  1176 => x"80ddc008",
  1177 => x"f80c881d",
  1178 => x"54807480",
  1179 => x"f52d7081",
  1180 => x"ff065558",
  1181 => x"5572752e",
  1182 => x"b6388114",
  1183 => x"80f52d53",
  1184 => x"72752eab",
  1185 => x"38748215",
  1186 => x"80f52d54",
  1187 => x"567280d3",
  1188 => x"2e098106",
  1189 => x"83388156",
  1190 => x"7280f332",
  1191 => x"70098105",
  1192 => x"70802578",
  1193 => x"07515153",
  1194 => x"72802e83",
  1195 => x"38a05580",
  1196 => x"7781ff06",
  1197 => x"54567280",
  1198 => x"c52e0981",
  1199 => x"06833881",
  1200 => x"567280e5",
  1201 => x"32700981",
  1202 => x"05708025",
  1203 => x"78075151",
  1204 => x"5372802e",
  1205 => x"a4388114",
  1206 => x"80f52d53",
  1207 => x"72b02e09",
  1208 => x"81068938",
  1209 => x"74828007",
  1210 => x"55a5f904",
  1211 => x"72b72e09",
  1212 => x"81068638",
  1213 => x"74848007",
  1214 => x"5580dbdc",
  1215 => x"08f9df06",
  1216 => x"750780db",
  1217 => x"dc0ca290",
  1218 => x"2d800be0",
  1219 => x"0c805186",
  1220 => x"da2d86c7",
  1221 => x"2d7a802e",
  1222 => x"883880d8",
  1223 => x"e051a6a5",
  1224 => x"0480da88",
  1225 => x"51b0ad2d",
  1226 => x"7a80dda0",
  1227 => x"0c02b405",
  1228 => x"0d0402f4",
  1229 => x"050d840b",
  1230 => x"ec0c810b",
  1231 => x"e00cadea",
  1232 => x"2da7c42d",
  1233 => x"81f92d83",
  1234 => x"52adcd2d",
  1235 => x"8151858d",
  1236 => x"2dff1252",
  1237 => x"718025f1",
  1238 => x"38840bec",
  1239 => x"0c80d790",
  1240 => x"5186a02d",
  1241 => x"80c2ab2d",
  1242 => x"80dda008",
  1243 => x"802ebe38",
  1244 => x"a3b45180",
  1245 => x"d5b12d80",
  1246 => x"d8e051b0",
  1247 => x"ad2dae8c",
  1248 => x"2da8ef2d",
  1249 => x"80dda008",
  1250 => x"81065271",
  1251 => x"802e8638",
  1252 => x"805194bf",
  1253 => x"2db0c02d",
  1254 => x"80dda008",
  1255 => x"52a2902d",
  1256 => x"86537183",
  1257 => x"38845372",
  1258 => x"ec0ca781",
  1259 => x"04800b80",
  1260 => x"dda00c02",
  1261 => x"8c050d04",
  1262 => x"71980c04",
  1263 => x"ffb00880",
  1264 => x"dda00c04",
  1265 => x"810bffb0",
  1266 => x"0c04800b",
  1267 => x"ffb00c04",
  1268 => x"02d8050d",
  1269 => x"ffb40887",
  1270 => x"ffff065a",
  1271 => x"81548070",
  1272 => x"80dbc808",
  1273 => x"80dbcc08",
  1274 => x"80dba45b",
  1275 => x"59575a58",
  1276 => x"79740675",
  1277 => x"75065252",
  1278 => x"71712e8d",
  1279 => x"38807781",
  1280 => x"8a2d7309",
  1281 => x"75067207",
  1282 => x"557680e0",
  1283 => x"2d7083ff",
  1284 => x"ff065351",
  1285 => x"7180e42e",
  1286 => x"098106a2",
  1287 => x"38747406",
  1288 => x"70777606",
  1289 => x"32700981",
  1290 => x"05707207",
  1291 => x"9f2a7b05",
  1292 => x"77097a06",
  1293 => x"74075a5b",
  1294 => x"535353a8",
  1295 => x"cc047180",
  1296 => x"e4268938",
  1297 => x"81115170",
  1298 => x"77818a2d",
  1299 => x"7310811a",
  1300 => x"8219595a",
  1301 => x"54907925",
  1302 => x"ff963875",
  1303 => x"80dbcc0c",
  1304 => x"7480dbc8",
  1305 => x"0c7780dd",
  1306 => x"a00c02a8",
  1307 => x"050d0402",
  1308 => x"d0050d80",
  1309 => x"5ca9ff04",
  1310 => x"80dda008",
  1311 => x"81f02e09",
  1312 => x"81068a38",
  1313 => x"810b80db",
  1314 => x"d40ca9ff",
  1315 => x"0480dda0",
  1316 => x"0881e02e",
  1317 => x"0981068a",
  1318 => x"38810b80",
  1319 => x"dbd80ca9",
  1320 => x"ff0480dd",
  1321 => x"a0085280",
  1322 => x"dbd80880",
  1323 => x"2e893880",
  1324 => x"dda00881",
  1325 => x"80055271",
  1326 => x"842c728f",
  1327 => x"06535380",
  1328 => x"dbd40880",
  1329 => x"2e9a3872",
  1330 => x"842980da",
  1331 => x"ac057213",
  1332 => x"81712b70",
  1333 => x"09730806",
  1334 => x"730c5153",
  1335 => x"53a9f304",
  1336 => x"72842980",
  1337 => x"daac0572",
  1338 => x"1383712b",
  1339 => x"72080772",
  1340 => x"0c535380",
  1341 => x"0b80dbd8",
  1342 => x"0c800b80",
  1343 => x"dbd40c80",
  1344 => x"ddc851ac",
  1345 => x"c02d80dd",
  1346 => x"a008ff24",
  1347 => x"feea38a7",
  1348 => x"d02d80dd",
  1349 => x"a008802e",
  1350 => x"81b03881",
  1351 => x"59800b80",
  1352 => x"dbd00880",
  1353 => x"dbcc0880",
  1354 => x"db805a5c",
  1355 => x"5c587a79",
  1356 => x"067a7a06",
  1357 => x"54527173",
  1358 => x"2e80f838",
  1359 => x"72098105",
  1360 => x"70740780",
  1361 => x"2580daec",
  1362 => x"1a80f52d",
  1363 => x"70842c71",
  1364 => x"8f065853",
  1365 => x"57575275",
  1366 => x"802ea338",
  1367 => x"71842980",
  1368 => x"daac0574",
  1369 => x"1583712b",
  1370 => x"72080772",
  1371 => x"0c545276",
  1372 => x"80e02d81",
  1373 => x"05527177",
  1374 => x"818a2dab",
  1375 => x"94047184",
  1376 => x"2980daac",
  1377 => x"05741581",
  1378 => x"712b7009",
  1379 => x"73080673",
  1380 => x"0c515353",
  1381 => x"74853270",
  1382 => x"09810570",
  1383 => x"80255151",
  1384 => x"5275802e",
  1385 => x"8e388170",
  1386 => x"73065353",
  1387 => x"71802e83",
  1388 => x"38725c78",
  1389 => x"10811982",
  1390 => x"19595959",
  1391 => x"907825fe",
  1392 => x"ed3880db",
  1393 => x"cc0880db",
  1394 => x"d00c7b80",
  1395 => x"dda00c02",
  1396 => x"b0050d04",
  1397 => x"02f8050d",
  1398 => x"80daac52",
  1399 => x"8f518072",
  1400 => x"70840554",
  1401 => x"0cff1151",
  1402 => x"708025f2",
  1403 => x"38028805",
  1404 => x"0d0402f0",
  1405 => x"050d7551",
  1406 => x"a7ca2d70",
  1407 => x"822cfc06",
  1408 => x"80daac11",
  1409 => x"72109e06",
  1410 => x"71087072",
  1411 => x"2a708306",
  1412 => x"82742b70",
  1413 => x"09740676",
  1414 => x"0c545156",
  1415 => x"57535153",
  1416 => x"a7c42d71",
  1417 => x"80dda00c",
  1418 => x"0290050d",
  1419 => x"0402fc05",
  1420 => x"0d725180",
  1421 => x"710c800b",
  1422 => x"84120c02",
  1423 => x"84050d04",
  1424 => x"02f0050d",
  1425 => x"75700884",
  1426 => x"12085353",
  1427 => x"53ff5471",
  1428 => x"712ea838",
  1429 => x"a7ca2d84",
  1430 => x"13087084",
  1431 => x"29148811",
  1432 => x"70087081",
  1433 => x"ff068418",
  1434 => x"08811187",
  1435 => x"06841a0c",
  1436 => x"53515551",
  1437 => x"5151a7c4",
  1438 => x"2d715473",
  1439 => x"80dda00c",
  1440 => x"0290050d",
  1441 => x"0402f805",
  1442 => x"0da7ca2d",
  1443 => x"e008708b",
  1444 => x"2a708106",
  1445 => x"51525270",
  1446 => x"802ea138",
  1447 => x"80ddc808",
  1448 => x"70842980",
  1449 => x"ddd00573",
  1450 => x"81ff0671",
  1451 => x"0c515180",
  1452 => x"ddc80881",
  1453 => x"11870680",
  1454 => x"ddc80c51",
  1455 => x"800b80dd",
  1456 => x"f00ca7bc",
  1457 => x"2da7c42d",
  1458 => x"0288050d",
  1459 => x"0402fc05",
  1460 => x"0da7ca2d",
  1461 => x"810b80dd",
  1462 => x"f00ca7c4",
  1463 => x"2d80ddf0",
  1464 => x"085170f9",
  1465 => x"38028405",
  1466 => x"0d0402fc",
  1467 => x"050d80dd",
  1468 => x"c851acad",
  1469 => x"2dabd42d",
  1470 => x"ad8551a7",
  1471 => x"b82d0284",
  1472 => x"050d0480",
  1473 => x"ddfc0880",
  1474 => x"dda00c04",
  1475 => x"02fc050d",
  1476 => x"810b80db",
  1477 => x"e00c8151",
  1478 => x"858d2d02",
  1479 => x"84050d04",
  1480 => x"02fc050d",
  1481 => x"aeaa04a8",
  1482 => x"ef2d80f6",
  1483 => x"51abf22d",
  1484 => x"80dda008",
  1485 => x"f23880da",
  1486 => x"51abf22d",
  1487 => x"80dda008",
  1488 => x"e63880dd",
  1489 => x"a00880db",
  1490 => x"e00c80dd",
  1491 => x"a0085185",
  1492 => x"8d2d0284",
  1493 => x"050d0402",
  1494 => x"ec050d76",
  1495 => x"54805287",
  1496 => x"0b881580",
  1497 => x"f52d5653",
  1498 => x"74722483",
  1499 => x"38a05372",
  1500 => x"5183842d",
  1501 => x"81128b15",
  1502 => x"80f52d54",
  1503 => x"52727225",
  1504 => x"de380294",
  1505 => x"050d0402",
  1506 => x"f0050d80",
  1507 => x"ddfc0854",
  1508 => x"81f92d80",
  1509 => x"0b80de80",
  1510 => x"0c730880",
  1511 => x"2e818938",
  1512 => x"820b80dd",
  1513 => x"b40c80de",
  1514 => x"80088f06",
  1515 => x"80ddb00c",
  1516 => x"73085271",
  1517 => x"832e9638",
  1518 => x"71832689",
  1519 => x"3871812e",
  1520 => x"b038b091",
  1521 => x"0471852e",
  1522 => x"a038b091",
  1523 => x"04881480",
  1524 => x"f52d8415",
  1525 => x"0880d7a8",
  1526 => x"53545286",
  1527 => x"a02d7184",
  1528 => x"29137008",
  1529 => x"5252b095",
  1530 => x"047351ae",
  1531 => x"d72db091",
  1532 => x"0480dbdc",
  1533 => x"08881508",
  1534 => x"2c708106",
  1535 => x"51527180",
  1536 => x"2e883880",
  1537 => x"d7ac51b0",
  1538 => x"8e0480d7",
  1539 => x"b05186a0",
  1540 => x"2d841408",
  1541 => x"5186a02d",
  1542 => x"80de8008",
  1543 => x"810580de",
  1544 => x"800c8c14",
  1545 => x"54af9904",
  1546 => x"0290050d",
  1547 => x"047180dd",
  1548 => x"fc0caf87",
  1549 => x"2d80de80",
  1550 => x"08ff0580",
  1551 => x"de840c04",
  1552 => x"02e8050d",
  1553 => x"80ddfc08",
  1554 => x"80de8808",
  1555 => x"575580f6",
  1556 => x"51abf22d",
  1557 => x"80dda008",
  1558 => x"812a7081",
  1559 => x"06515271",
  1560 => x"802ea438",
  1561 => x"b0ea04a8",
  1562 => x"ef2d80f6",
  1563 => x"51abf22d",
  1564 => x"80dda008",
  1565 => x"f23880db",
  1566 => x"e0088132",
  1567 => x"7080dbe0",
  1568 => x"0c705252",
  1569 => x"858d2d80",
  1570 => x"0b80ddf4",
  1571 => x"0c800b80",
  1572 => x"ddf80c80",
  1573 => x"dbe00883",
  1574 => x"8d3880da",
  1575 => x"51abf22d",
  1576 => x"80dda008",
  1577 => x"802e8c38",
  1578 => x"80ddf408",
  1579 => x"81800780",
  1580 => x"ddf40c80",
  1581 => x"d951abf2",
  1582 => x"2d80dda0",
  1583 => x"08802e8c",
  1584 => x"3880ddf4",
  1585 => x"0880c007",
  1586 => x"80ddf40c",
  1587 => x"819451ab",
  1588 => x"f22d80dd",
  1589 => x"a008802e",
  1590 => x"8b3880dd",
  1591 => x"f4089007",
  1592 => x"80ddf40c",
  1593 => x"819151ab",
  1594 => x"f22d80dd",
  1595 => x"a008802e",
  1596 => x"8b3880dd",
  1597 => x"f408a007",
  1598 => x"80ddf40c",
  1599 => x"81f551ab",
  1600 => x"f22d80dd",
  1601 => x"a008802e",
  1602 => x"8b3880dd",
  1603 => x"f4088107",
  1604 => x"80ddf40c",
  1605 => x"81f251ab",
  1606 => x"f22d80dd",
  1607 => x"a008802e",
  1608 => x"8b3880dd",
  1609 => x"f4088207",
  1610 => x"80ddf40c",
  1611 => x"81eb51ab",
  1612 => x"f22d80dd",
  1613 => x"a008802e",
  1614 => x"8b3880dd",
  1615 => x"f4088407",
  1616 => x"80ddf40c",
  1617 => x"81f451ab",
  1618 => x"f22d80dd",
  1619 => x"a008802e",
  1620 => x"8b3880dd",
  1621 => x"f4088807",
  1622 => x"80ddf40c",
  1623 => x"80d851ab",
  1624 => x"f22d80dd",
  1625 => x"a008802e",
  1626 => x"8c3880dd",
  1627 => x"f8088180",
  1628 => x"0780ddf8",
  1629 => x"0c9251ab",
  1630 => x"f22d80dd",
  1631 => x"a008802e",
  1632 => x"8c3880dd",
  1633 => x"f80880c0",
  1634 => x"0780ddf8",
  1635 => x"0c9451ab",
  1636 => x"f22d80dd",
  1637 => x"a008802e",
  1638 => x"8b3880dd",
  1639 => x"f8089007",
  1640 => x"80ddf80c",
  1641 => x"9151abf2",
  1642 => x"2d80dda0",
  1643 => x"08802e8b",
  1644 => x"3880ddf8",
  1645 => x"08a00780",
  1646 => x"ddf80c9d",
  1647 => x"51abf22d",
  1648 => x"80dda008",
  1649 => x"802e8b38",
  1650 => x"80ddf808",
  1651 => x"810780dd",
  1652 => x"f80c9b51",
  1653 => x"abf22d80",
  1654 => x"dda00880",
  1655 => x"2e8b3880",
  1656 => x"ddf80882",
  1657 => x"0780ddf8",
  1658 => x"0c9c51ab",
  1659 => x"f22d80dd",
  1660 => x"a008802e",
  1661 => x"8b3880dd",
  1662 => x"f8088407",
  1663 => x"80ddf80c",
  1664 => x"a351abf2",
  1665 => x"2d80dda0",
  1666 => x"08802e8b",
  1667 => x"3880ddf8",
  1668 => x"08880780",
  1669 => x"ddf80c81",
  1670 => x"fd51abf2",
  1671 => x"2d81fa51",
  1672 => x"abf22db9",
  1673 => x"fb0481f5",
  1674 => x"51abf22d",
  1675 => x"80dda008",
  1676 => x"812a7081",
  1677 => x"06515271",
  1678 => x"802eb338",
  1679 => x"80de8408",
  1680 => x"5271802e",
  1681 => x"8a38ff12",
  1682 => x"80de840c",
  1683 => x"b4ee0480",
  1684 => x"de800810",
  1685 => x"80de8008",
  1686 => x"05708429",
  1687 => x"16515288",
  1688 => x"1208802e",
  1689 => x"8938ff51",
  1690 => x"88120852",
  1691 => x"712d81f2",
  1692 => x"51abf22d",
  1693 => x"80dda008",
  1694 => x"812a7081",
  1695 => x"06515271",
  1696 => x"802eb438",
  1697 => x"80de8008",
  1698 => x"ff1180de",
  1699 => x"84085653",
  1700 => x"53737225",
  1701 => x"8a388114",
  1702 => x"80de840c",
  1703 => x"b5b70472",
  1704 => x"10137084",
  1705 => x"29165152",
  1706 => x"88120880",
  1707 => x"2e8938fe",
  1708 => x"51881208",
  1709 => x"52712d81",
  1710 => x"fd51abf2",
  1711 => x"2d80dda0",
  1712 => x"08812a70",
  1713 => x"81065152",
  1714 => x"71802eb1",
  1715 => x"3880de84",
  1716 => x"08802e8a",
  1717 => x"38800b80",
  1718 => x"de840cb5",
  1719 => x"fd0480de",
  1720 => x"80081080",
  1721 => x"de800805",
  1722 => x"70842916",
  1723 => x"51528812",
  1724 => x"08802e89",
  1725 => x"38fd5188",
  1726 => x"12085271",
  1727 => x"2d81fa51",
  1728 => x"abf22d80",
  1729 => x"dda00881",
  1730 => x"2a708106",
  1731 => x"51527180",
  1732 => x"2eb13880",
  1733 => x"de8008ff",
  1734 => x"11545280",
  1735 => x"de840873",
  1736 => x"25893872",
  1737 => x"80de840c",
  1738 => x"b6c30471",
  1739 => x"10127084",
  1740 => x"29165152",
  1741 => x"88120880",
  1742 => x"2e8938fc",
  1743 => x"51881208",
  1744 => x"52712d80",
  1745 => x"de840870",
  1746 => x"53547380",
  1747 => x"2e8a388c",
  1748 => x"15ff1555",
  1749 => x"55b6ca04",
  1750 => x"820b80dd",
  1751 => x"b40c718f",
  1752 => x"0680ddb0",
  1753 => x"0c81eb51",
  1754 => x"abf22d80",
  1755 => x"dda00881",
  1756 => x"2a708106",
  1757 => x"51527180",
  1758 => x"2ead3874",
  1759 => x"08852e09",
  1760 => x"8106a438",
  1761 => x"881580f5",
  1762 => x"2dff0552",
  1763 => x"71881681",
  1764 => x"b72d7198",
  1765 => x"2b527180",
  1766 => x"25883880",
  1767 => x"0b881681",
  1768 => x"b72d7451",
  1769 => x"aed72d81",
  1770 => x"f451abf2",
  1771 => x"2d80dda0",
  1772 => x"08812a70",
  1773 => x"81065152",
  1774 => x"71802eb3",
  1775 => x"38740885",
  1776 => x"2e098106",
  1777 => x"aa388815",
  1778 => x"80f52d81",
  1779 => x"05527188",
  1780 => x"1681b72d",
  1781 => x"7181ff06",
  1782 => x"8b1680f5",
  1783 => x"2d545272",
  1784 => x"72278738",
  1785 => x"72881681",
  1786 => x"b72d7451",
  1787 => x"aed72d80",
  1788 => x"da51abf2",
  1789 => x"2d80dda0",
  1790 => x"08812a70",
  1791 => x"81065152",
  1792 => x"71802e81",
  1793 => x"ad3880dd",
  1794 => x"fc0880de",
  1795 => x"84085553",
  1796 => x"73802e8a",
  1797 => x"388c13ff",
  1798 => x"155553b8",
  1799 => x"90047208",
  1800 => x"5271822e",
  1801 => x"a6387182",
  1802 => x"26893871",
  1803 => x"812eaa38",
  1804 => x"b9b20471",
  1805 => x"832eb438",
  1806 => x"71842e09",
  1807 => x"810680f2",
  1808 => x"38881308",
  1809 => x"51b0ad2d",
  1810 => x"b9b20480",
  1811 => x"de840851",
  1812 => x"88130852",
  1813 => x"712db9b2",
  1814 => x"04810b88",
  1815 => x"14082b80",
  1816 => x"dbdc0832",
  1817 => x"80dbdc0c",
  1818 => x"b9860488",
  1819 => x"1380f52d",
  1820 => x"81058b14",
  1821 => x"80f52d53",
  1822 => x"54717424",
  1823 => x"83388054",
  1824 => x"73881481",
  1825 => x"b72daf87",
  1826 => x"2db9b204",
  1827 => x"7508802e",
  1828 => x"a4387508",
  1829 => x"51abf22d",
  1830 => x"80dda008",
  1831 => x"81065271",
  1832 => x"802e8c38",
  1833 => x"80de8408",
  1834 => x"51841608",
  1835 => x"52712d88",
  1836 => x"165675d8",
  1837 => x"38805480",
  1838 => x"0b80ddb4",
  1839 => x"0c738f06",
  1840 => x"80ddb00c",
  1841 => x"a0527380",
  1842 => x"de84082e",
  1843 => x"09810699",
  1844 => x"3880de80",
  1845 => x"08ff0574",
  1846 => x"32700981",
  1847 => x"05707207",
  1848 => x"9f2a9171",
  1849 => x"31515153",
  1850 => x"53715183",
  1851 => x"842d8114",
  1852 => x"548e7425",
  1853 => x"c23880db",
  1854 => x"e0085271",
  1855 => x"80dda00c",
  1856 => x"0298050d",
  1857 => x"0402f405",
  1858 => x"0dd45281",
  1859 => x"ff720c71",
  1860 => x"085381ff",
  1861 => x"720c7288",
  1862 => x"2b83fe80",
  1863 => x"06720870",
  1864 => x"81ff0651",
  1865 => x"525381ff",
  1866 => x"720c7271",
  1867 => x"07882b72",
  1868 => x"087081ff",
  1869 => x"06515253",
  1870 => x"81ff720c",
  1871 => x"72710788",
  1872 => x"2b720870",
  1873 => x"81ff0672",
  1874 => x"0780dda0",
  1875 => x"0c525302",
  1876 => x"8c050d04",
  1877 => x"02f4050d",
  1878 => x"74767181",
  1879 => x"ff06d40c",
  1880 => x"535380de",
  1881 => x"8c088538",
  1882 => x"71892b52",
  1883 => x"71982ad4",
  1884 => x"0c71902a",
  1885 => x"7081ff06",
  1886 => x"d40c5171",
  1887 => x"882a7081",
  1888 => x"ff06d40c",
  1889 => x"517181ff",
  1890 => x"06d40c72",
  1891 => x"902a7081",
  1892 => x"ff06d40c",
  1893 => x"51d40870",
  1894 => x"81ff0651",
  1895 => x"5182b8bf",
  1896 => x"527081ff",
  1897 => x"2e098106",
  1898 => x"943881ff",
  1899 => x"0bd40cd4",
  1900 => x"087081ff",
  1901 => x"06ff1454",
  1902 => x"515171e5",
  1903 => x"387080dd",
  1904 => x"a00c028c",
  1905 => x"050d0402",
  1906 => x"fc050d81",
  1907 => x"c75181ff",
  1908 => x"0bd40cff",
  1909 => x"11517080",
  1910 => x"25f43802",
  1911 => x"84050d04",
  1912 => x"02f4050d",
  1913 => x"81ff0bd4",
  1914 => x"0c935380",
  1915 => x"5287fc80",
  1916 => x"c151bad4",
  1917 => x"2d80dda0",
  1918 => x"088b3881",
  1919 => x"ff0bd40c",
  1920 => x"8153bc8e",
  1921 => x"04bbc72d",
  1922 => x"ff135372",
  1923 => x"de387280",
  1924 => x"dda00c02",
  1925 => x"8c050d04",
  1926 => x"02ec050d",
  1927 => x"810b80de",
  1928 => x"8c0c8454",
  1929 => x"d008708f",
  1930 => x"2a708106",
  1931 => x"51515372",
  1932 => x"f33872d0",
  1933 => x"0cbbc72d",
  1934 => x"80d7b451",
  1935 => x"86a02dd0",
  1936 => x"08708f2a",
  1937 => x"70810651",
  1938 => x"515372f3",
  1939 => x"38810bd0",
  1940 => x"0cb15380",
  1941 => x"5284d480",
  1942 => x"c051bad4",
  1943 => x"2d80dda0",
  1944 => x"08812e93",
  1945 => x"3872822e",
  1946 => x"bf38ff13",
  1947 => x"5372e438",
  1948 => x"ff145473",
  1949 => x"ffae38bb",
  1950 => x"c72d83aa",
  1951 => x"52849c80",
  1952 => x"c851bad4",
  1953 => x"2d80dda0",
  1954 => x"08812e09",
  1955 => x"81069338",
  1956 => x"ba852d80",
  1957 => x"dda00883",
  1958 => x"ffff0653",
  1959 => x"7283aa2e",
  1960 => x"9f38bbe0",
  1961 => x"2dbdbb04",
  1962 => x"80d7c051",
  1963 => x"86a02d80",
  1964 => x"53bf9004",
  1965 => x"80d7d851",
  1966 => x"86a02d80",
  1967 => x"54bee104",
  1968 => x"81ff0bd4",
  1969 => x"0cb154bb",
  1970 => x"c72d8fcf",
  1971 => x"53805287",
  1972 => x"fc80f751",
  1973 => x"bad42d80",
  1974 => x"dda00855",
  1975 => x"80dda008",
  1976 => x"812e0981",
  1977 => x"069c3881",
  1978 => x"ff0bd40c",
  1979 => x"820a5284",
  1980 => x"9c80e951",
  1981 => x"bad42d80",
  1982 => x"dda00880",
  1983 => x"2e8d38bb",
  1984 => x"c72dff13",
  1985 => x"5372c638",
  1986 => x"bed40481",
  1987 => x"ff0bd40c",
  1988 => x"80dda008",
  1989 => x"5287fc80",
  1990 => x"fa51bad4",
  1991 => x"2d80dda0",
  1992 => x"08b23881",
  1993 => x"ff0bd40c",
  1994 => x"d4085381",
  1995 => x"ff0bd40c",
  1996 => x"81ff0bd4",
  1997 => x"0c81ff0b",
  1998 => x"d40c81ff",
  1999 => x"0bd40c72",
  2000 => x"862a7081",
  2001 => x"06765651",
  2002 => x"53729638",
  2003 => x"80dda008",
  2004 => x"54bee104",
  2005 => x"73822efe",
  2006 => x"db38ff14",
  2007 => x"5473fee7",
  2008 => x"387380de",
  2009 => x"8c0c738b",
  2010 => x"38815287",
  2011 => x"fc80d051",
  2012 => x"bad42d81",
  2013 => x"ff0bd40c",
  2014 => x"d008708f",
  2015 => x"2a708106",
  2016 => x"51515372",
  2017 => x"f33872d0",
  2018 => x"0c81ff0b",
  2019 => x"d40c8153",
  2020 => x"7280dda0",
  2021 => x"0c029405",
  2022 => x"0d0402e8",
  2023 => x"050d7855",
  2024 => x"805681ff",
  2025 => x"0bd40cd0",
  2026 => x"08708f2a",
  2027 => x"70810651",
  2028 => x"515372f3",
  2029 => x"3882810b",
  2030 => x"d00c81ff",
  2031 => x"0bd40c77",
  2032 => x"5287fc80",
  2033 => x"d151bad4",
  2034 => x"2d80dbc6",
  2035 => x"df5480dd",
  2036 => x"a008802e",
  2037 => x"8c3880d7",
  2038 => x"f85186a0",
  2039 => x"2d80c0b6",
  2040 => x"0481ff0b",
  2041 => x"d40cd408",
  2042 => x"7081ff06",
  2043 => x"51537281",
  2044 => x"fe2e0981",
  2045 => x"069f3880",
  2046 => x"ff53ba85",
  2047 => x"2d80dda0",
  2048 => x"08757084",
  2049 => x"05570cff",
  2050 => x"13537280",
  2051 => x"25ec3881",
  2052 => x"5680c09b",
  2053 => x"04ff1454",
  2054 => x"73c73881",
  2055 => x"ff0bd40c",
  2056 => x"81ff0bd4",
  2057 => x"0cd00870",
  2058 => x"8f2a7081",
  2059 => x"06515153",
  2060 => x"72f33872",
  2061 => x"d00c7580",
  2062 => x"dda00c02",
  2063 => x"98050d04",
  2064 => x"02e8050d",
  2065 => x"77797b58",
  2066 => x"55558053",
  2067 => x"727625a5",
  2068 => x"38747081",
  2069 => x"055680f5",
  2070 => x"2d747081",
  2071 => x"055680f5",
  2072 => x"2d525271",
  2073 => x"712e8738",
  2074 => x"815180c0",
  2075 => x"f7048113",
  2076 => x"5380c0cc",
  2077 => x"04805170",
  2078 => x"80dda00c",
  2079 => x"0298050d",
  2080 => x"0402ec05",
  2081 => x"0d765574",
  2082 => x"802e80c4",
  2083 => x"389a1580",
  2084 => x"e02d5180",
  2085 => x"cfb52d80",
  2086 => x"dda00880",
  2087 => x"dda00880",
  2088 => x"e4c00c80",
  2089 => x"dda00854",
  2090 => x"5480e49c",
  2091 => x"08802e9b",
  2092 => x"38941580",
  2093 => x"e02d5180",
  2094 => x"cfb52d80",
  2095 => x"dda00890",
  2096 => x"2b83fff0",
  2097 => x"0a067075",
  2098 => x"07515372",
  2099 => x"80e4c00c",
  2100 => x"80e4c008",
  2101 => x"5372802e",
  2102 => x"9e3880e4",
  2103 => x"9408fe14",
  2104 => x"712980e4",
  2105 => x"a8080580",
  2106 => x"e4c40c70",
  2107 => x"842b80e4",
  2108 => x"a00c5480",
  2109 => x"c2a60480",
  2110 => x"e4ac0880",
  2111 => x"e4c00c80",
  2112 => x"e4b00880",
  2113 => x"e4c40c80",
  2114 => x"e49c0880",
  2115 => x"2e8c3880",
  2116 => x"e4940884",
  2117 => x"2b5380c2",
  2118 => x"a10480e4",
  2119 => x"b408842b",
  2120 => x"537280e4",
  2121 => x"a00c0294",
  2122 => x"050d0402",
  2123 => x"d8050d80",
  2124 => x"0b80e49c",
  2125 => x"0c8454bc",
  2126 => x"982d80dd",
  2127 => x"a008802e",
  2128 => x"983880de",
  2129 => x"90528051",
  2130 => x"bf9a2d80",
  2131 => x"dda00880",
  2132 => x"2e8738fe",
  2133 => x"5480c2e1",
  2134 => x"04ff1454",
  2135 => x"738024d7",
  2136 => x"38738e38",
  2137 => x"80d88851",
  2138 => x"86a02d73",
  2139 => x"5580c8c4",
  2140 => x"04805681",
  2141 => x"0b80e4c8",
  2142 => x"0c885380",
  2143 => x"d89c5280",
  2144 => x"dec65180",
  2145 => x"c0c02d80",
  2146 => x"dda00876",
  2147 => x"2e098106",
  2148 => x"893880dd",
  2149 => x"a00880e4",
  2150 => x"c80c8853",
  2151 => x"80d8a852",
  2152 => x"80dee251",
  2153 => x"80c0c02d",
  2154 => x"80dda008",
  2155 => x"893880dd",
  2156 => x"a00880e4",
  2157 => x"c80c80e4",
  2158 => x"c808802e",
  2159 => x"81843880",
  2160 => x"e1d60b80",
  2161 => x"f52d80e1",
  2162 => x"d70b80f5",
  2163 => x"2d71982b",
  2164 => x"71902b07",
  2165 => x"80e1d80b",
  2166 => x"80f52d70",
  2167 => x"882b7207",
  2168 => x"80e1d90b",
  2169 => x"80f52d71",
  2170 => x"0780e28e",
  2171 => x"0b80f52d",
  2172 => x"80e28f0b",
  2173 => x"80f52d71",
  2174 => x"882b0753",
  2175 => x"5f54525a",
  2176 => x"56575573",
  2177 => x"81abaa2e",
  2178 => x"09810690",
  2179 => x"38755180",
  2180 => x"cf842d80",
  2181 => x"dda00856",
  2182 => x"80c4ab04",
  2183 => x"7382d4d5",
  2184 => x"2e893880",
  2185 => x"d8b45180",
  2186 => x"c4fa0480",
  2187 => x"de905275",
  2188 => x"51bf9a2d",
  2189 => x"80dda008",
  2190 => x"5580dda0",
  2191 => x"08802e84",
  2192 => x"83388853",
  2193 => x"80d8a852",
  2194 => x"80dee251",
  2195 => x"80c0c02d",
  2196 => x"80dda008",
  2197 => x"8b38810b",
  2198 => x"80e49c0c",
  2199 => x"80c58104",
  2200 => x"885380d8",
  2201 => x"9c5280de",
  2202 => x"c65180c0",
  2203 => x"c02d80dd",
  2204 => x"a008802e",
  2205 => x"8c3880d8",
  2206 => x"c85186a0",
  2207 => x"2d80c5e0",
  2208 => x"0480e28e",
  2209 => x"0b80f52d",
  2210 => x"547380d5",
  2211 => x"2e098106",
  2212 => x"80ce3880",
  2213 => x"e28f0b80",
  2214 => x"f52d5473",
  2215 => x"81aa2e09",
  2216 => x"8106bd38",
  2217 => x"800b80de",
  2218 => x"900b80f5",
  2219 => x"2d565474",
  2220 => x"81e92e83",
  2221 => x"38815474",
  2222 => x"81eb2e8c",
  2223 => x"38805573",
  2224 => x"752e0981",
  2225 => x"0682fd38",
  2226 => x"80de9b0b",
  2227 => x"80f52d55",
  2228 => x"748e3880",
  2229 => x"de9c0b80",
  2230 => x"f52d5473",
  2231 => x"822e8738",
  2232 => x"805580c8",
  2233 => x"c40480de",
  2234 => x"9d0b80f5",
  2235 => x"2d7080e4",
  2236 => x"940cff05",
  2237 => x"80e4980c",
  2238 => x"80de9e0b",
  2239 => x"80f52d80",
  2240 => x"de9f0b80",
  2241 => x"f52d5876",
  2242 => x"05778280",
  2243 => x"29057080",
  2244 => x"e4a40c80",
  2245 => x"dea00b80",
  2246 => x"f52d7080",
  2247 => x"e4b80c80",
  2248 => x"e49c0859",
  2249 => x"57587680",
  2250 => x"2e81b938",
  2251 => x"885380d8",
  2252 => x"a85280de",
  2253 => x"e25180c0",
  2254 => x"c02d80dd",
  2255 => x"a0088284",
  2256 => x"3880e494",
  2257 => x"0870842b",
  2258 => x"80e4a00c",
  2259 => x"7080e4b4",
  2260 => x"0c80deb5",
  2261 => x"0b80f52d",
  2262 => x"80deb40b",
  2263 => x"80f52d71",
  2264 => x"82802905",
  2265 => x"80deb60b",
  2266 => x"80f52d70",
  2267 => x"84808029",
  2268 => x"1280deb7",
  2269 => x"0b80f52d",
  2270 => x"7081800a",
  2271 => x"29127080",
  2272 => x"e4bc0c80",
  2273 => x"e4b80871",
  2274 => x"2980e4a4",
  2275 => x"08057080",
  2276 => x"e4a80c80",
  2277 => x"debd0b80",
  2278 => x"f52d80de",
  2279 => x"bc0b80f5",
  2280 => x"2d718280",
  2281 => x"290580de",
  2282 => x"be0b80f5",
  2283 => x"2d708480",
  2284 => x"80291280",
  2285 => x"debf0b80",
  2286 => x"f52d7098",
  2287 => x"2b81f00a",
  2288 => x"06720570",
  2289 => x"80e4ac0c",
  2290 => x"fe117e29",
  2291 => x"770580e4",
  2292 => x"b00c5259",
  2293 => x"5243545e",
  2294 => x"51525952",
  2295 => x"5d575957",
  2296 => x"80c8bc04",
  2297 => x"80dea20b",
  2298 => x"80f52d80",
  2299 => x"dea10b80",
  2300 => x"f52d7182",
  2301 => x"80290570",
  2302 => x"80e4a00c",
  2303 => x"70a02983",
  2304 => x"ff057089",
  2305 => x"2a7080e4",
  2306 => x"b40c80de",
  2307 => x"a70b80f5",
  2308 => x"2d80dea6",
  2309 => x"0b80f52d",
  2310 => x"71828029",
  2311 => x"057080e4",
  2312 => x"bc0c7b71",
  2313 => x"291e7080",
  2314 => x"e4b00c7d",
  2315 => x"80e4ac0c",
  2316 => x"730580e4",
  2317 => x"a80c555e",
  2318 => x"51515555",
  2319 => x"805180c1",
  2320 => x"812d8155",
  2321 => x"7480dda0",
  2322 => x"0c02a805",
  2323 => x"0d0402ec",
  2324 => x"050d7670",
  2325 => x"872c7180",
  2326 => x"ff065556",
  2327 => x"5480e49c",
  2328 => x"088a3873",
  2329 => x"882c7481",
  2330 => x"ff065455",
  2331 => x"80de9052",
  2332 => x"80e4a408",
  2333 => x"1551bf9a",
  2334 => x"2d80dda0",
  2335 => x"085480dd",
  2336 => x"a008802e",
  2337 => x"bb3880e4",
  2338 => x"9c08802e",
  2339 => x"9c387284",
  2340 => x"2980de90",
  2341 => x"05700852",
  2342 => x"5380cf84",
  2343 => x"2d80dda0",
  2344 => x"08f00a06",
  2345 => x"5380c9be",
  2346 => x"04721080",
  2347 => x"de900570",
  2348 => x"80e02d52",
  2349 => x"5380cfb5",
  2350 => x"2d80dda0",
  2351 => x"08537254",
  2352 => x"7380dda0",
  2353 => x"0c029405",
  2354 => x"0d0402e0",
  2355 => x"050d7970",
  2356 => x"842c80e4",
  2357 => x"c4080571",
  2358 => x"8f065255",
  2359 => x"53728a38",
  2360 => x"80de9052",
  2361 => x"7351bf9a",
  2362 => x"2d72a029",
  2363 => x"80de9005",
  2364 => x"54807480",
  2365 => x"f52d5653",
  2366 => x"74732e83",
  2367 => x"38815374",
  2368 => x"81e52e81",
  2369 => x"f5388170",
  2370 => x"74065458",
  2371 => x"72802e81",
  2372 => x"e9388b14",
  2373 => x"80f52d70",
  2374 => x"832a7906",
  2375 => x"5856769c",
  2376 => x"3880dbe4",
  2377 => x"08537289",
  2378 => x"387280e2",
  2379 => x"900b81b7",
  2380 => x"2d7680db",
  2381 => x"e40c7353",
  2382 => x"80cbfc04",
  2383 => x"758f2e09",
  2384 => x"810681b6",
  2385 => x"38749f06",
  2386 => x"8d2980e2",
  2387 => x"83115153",
  2388 => x"811480f5",
  2389 => x"2d737081",
  2390 => x"055581b7",
  2391 => x"2d831480",
  2392 => x"f52d7370",
  2393 => x"81055581",
  2394 => x"b72d8514",
  2395 => x"80f52d73",
  2396 => x"70810555",
  2397 => x"81b72d87",
  2398 => x"1480f52d",
  2399 => x"73708105",
  2400 => x"5581b72d",
  2401 => x"891480f5",
  2402 => x"2d737081",
  2403 => x"055581b7",
  2404 => x"2d8e1480",
  2405 => x"f52d7370",
  2406 => x"81055581",
  2407 => x"b72d9014",
  2408 => x"80f52d73",
  2409 => x"70810555",
  2410 => x"81b72d92",
  2411 => x"1480f52d",
  2412 => x"73708105",
  2413 => x"5581b72d",
  2414 => x"941480f5",
  2415 => x"2d737081",
  2416 => x"055581b7",
  2417 => x"2d961480",
  2418 => x"f52d7370",
  2419 => x"81055581",
  2420 => x"b72d9814",
  2421 => x"80f52d73",
  2422 => x"70810555",
  2423 => x"81b72d9c",
  2424 => x"1480f52d",
  2425 => x"73708105",
  2426 => x"5581b72d",
  2427 => x"9e1480f5",
  2428 => x"2d7381b7",
  2429 => x"2d7780db",
  2430 => x"e40c8053",
  2431 => x"7280dda0",
  2432 => x"0c02a005",
  2433 => x"0d0402cc",
  2434 => x"050d7e60",
  2435 => x"5e5a800b",
  2436 => x"80e4c008",
  2437 => x"80e4c408",
  2438 => x"595c5680",
  2439 => x"5880e4a0",
  2440 => x"08782e81",
  2441 => x"bd38778f",
  2442 => x"06a01757",
  2443 => x"54739138",
  2444 => x"80de9052",
  2445 => x"76518117",
  2446 => x"57bf9a2d",
  2447 => x"80de9056",
  2448 => x"807680f5",
  2449 => x"2d565474",
  2450 => x"742e8338",
  2451 => x"81547481",
  2452 => x"e52e8182",
  2453 => x"38817075",
  2454 => x"06555c73",
  2455 => x"802e80f6",
  2456 => x"388b1680",
  2457 => x"f52d9806",
  2458 => x"597880ea",
  2459 => x"388b537c",
  2460 => x"52755180",
  2461 => x"c0c02d80",
  2462 => x"dda00880",
  2463 => x"d9389c16",
  2464 => x"085180cf",
  2465 => x"842d80dd",
  2466 => x"a008841b",
  2467 => x"0c9a1680",
  2468 => x"e02d5180",
  2469 => x"cfb52d80",
  2470 => x"dda00880",
  2471 => x"dda00888",
  2472 => x"1c0c80dd",
  2473 => x"a0085555",
  2474 => x"80e49c08",
  2475 => x"802e9a38",
  2476 => x"941680e0",
  2477 => x"2d5180cf",
  2478 => x"b52d80dd",
  2479 => x"a008902b",
  2480 => x"83fff00a",
  2481 => x"06701651",
  2482 => x"5473881b",
  2483 => x"0c787a0c",
  2484 => x"7b5480ce",
  2485 => x"a0048118",
  2486 => x"5880e4a0",
  2487 => x"087826fe",
  2488 => x"c53880e4",
  2489 => x"9c08802e",
  2490 => x"b5387a51",
  2491 => x"80c8ce2d",
  2492 => x"80dda008",
  2493 => x"80dda008",
  2494 => x"80ffffff",
  2495 => x"f806555b",
  2496 => x"7380ffff",
  2497 => x"fff82e96",
  2498 => x"3880dda0",
  2499 => x"08fe0580",
  2500 => x"e4940829",
  2501 => x"80e4a808",
  2502 => x"055780cc",
  2503 => x"9b048054",
  2504 => x"7380dda0",
  2505 => x"0c02b405",
  2506 => x"0d0402f4",
  2507 => x"050d7470",
  2508 => x"08810571",
  2509 => x"0c700880",
  2510 => x"e4980806",
  2511 => x"53537190",
  2512 => x"38881308",
  2513 => x"5180c8ce",
  2514 => x"2d80dda0",
  2515 => x"0888140c",
  2516 => x"810b80dd",
  2517 => x"a00c028c",
  2518 => x"050d0402",
  2519 => x"f0050d75",
  2520 => x"881108fe",
  2521 => x"0580e494",
  2522 => x"082980e4",
  2523 => x"a8081172",
  2524 => x"0880e498",
  2525 => x"08060579",
  2526 => x"55535454",
  2527 => x"bf9a2d02",
  2528 => x"90050d04",
  2529 => x"02f4050d",
  2530 => x"7470882a",
  2531 => x"83fe8006",
  2532 => x"7072982a",
  2533 => x"0772882b",
  2534 => x"87fc8080",
  2535 => x"0673982b",
  2536 => x"81f00a06",
  2537 => x"71730707",
  2538 => x"80dda00c",
  2539 => x"56515351",
  2540 => x"028c050d",
  2541 => x"0402f805",
  2542 => x"0d028e05",
  2543 => x"80f52d74",
  2544 => x"882b0770",
  2545 => x"83ffff06",
  2546 => x"80dda00c",
  2547 => x"51028805",
  2548 => x"0d0402f4",
  2549 => x"050d7476",
  2550 => x"78535452",
  2551 => x"80712597",
  2552 => x"38727081",
  2553 => x"055480f5",
  2554 => x"2d727081",
  2555 => x"055481b7",
  2556 => x"2dff1151",
  2557 => x"70eb3880",
  2558 => x"7281b72d",
  2559 => x"028c050d",
  2560 => x"0402e805",
  2561 => x"0d775680",
  2562 => x"70565473",
  2563 => x"7624b738",
  2564 => x"80e4a008",
  2565 => x"742eaf38",
  2566 => x"735180c9",
  2567 => x"ca2d80dd",
  2568 => x"a00880dd",
  2569 => x"a0080981",
  2570 => x"057080dd",
  2571 => x"a008079f",
  2572 => x"2a770581",
  2573 => x"17575753",
  2574 => x"53747624",
  2575 => x"893880e4",
  2576 => x"a0087426",
  2577 => x"d3387280",
  2578 => x"dda00c02",
  2579 => x"98050d04",
  2580 => x"02f0050d",
  2581 => x"80dd9c08",
  2582 => x"165180d0",
  2583 => x"812d80dd",
  2584 => x"a008802e",
  2585 => x"a0388b53",
  2586 => x"80dda008",
  2587 => x"5280e290",
  2588 => x"5180cfd2",
  2589 => x"2d80e4cc",
  2590 => x"08547380",
  2591 => x"2e873880",
  2592 => x"e2905173",
  2593 => x"2d029005",
  2594 => x"0d0402dc",
  2595 => x"050d8070",
  2596 => x"5a557480",
  2597 => x"dd9c0825",
  2598 => x"b53880e4",
  2599 => x"a008752e",
  2600 => x"ad387851",
  2601 => x"80c9ca2d",
  2602 => x"80dda008",
  2603 => x"09810570",
  2604 => x"80dda008",
  2605 => x"079f2a76",
  2606 => x"05811b5b",
  2607 => x"56547480",
  2608 => x"dd9c0825",
  2609 => x"893880e4",
  2610 => x"a0087926",
  2611 => x"d5388055",
  2612 => x"7880e4a0",
  2613 => x"082781e4",
  2614 => x"38785180",
  2615 => x"c9ca2d80",
  2616 => x"dda00880",
  2617 => x"2e81b438",
  2618 => x"80dda008",
  2619 => x"8b0580f5",
  2620 => x"2d70842a",
  2621 => x"70810677",
  2622 => x"1078842b",
  2623 => x"80e2900b",
  2624 => x"80f52d5c",
  2625 => x"5c535155",
  2626 => x"5673802e",
  2627 => x"80ce3874",
  2628 => x"16822b80",
  2629 => x"d3e00b80",
  2630 => x"dbf0120c",
  2631 => x"54777531",
  2632 => x"1080e4d0",
  2633 => x"11555690",
  2634 => x"74708105",
  2635 => x"5681b72d",
  2636 => x"a07481b7",
  2637 => x"2d7681ff",
  2638 => x"06811658",
  2639 => x"5473802e",
  2640 => x"8b389c53",
  2641 => x"80e29052",
  2642 => x"80d2d304",
  2643 => x"8b5380dd",
  2644 => x"a0085280",
  2645 => x"e4d21651",
  2646 => x"80d39104",
  2647 => x"7416822b",
  2648 => x"80d0d00b",
  2649 => x"80dbf012",
  2650 => x"0c547681",
  2651 => x"ff068116",
  2652 => x"58547380",
  2653 => x"2e8b389c",
  2654 => x"5380e290",
  2655 => x"5280d388",
  2656 => x"048b5380",
  2657 => x"dda00852",
  2658 => x"77753110",
  2659 => x"80e4d005",
  2660 => x"51765580",
  2661 => x"cfd22d80",
  2662 => x"d3b00474",
  2663 => x"90297531",
  2664 => x"701080e4",
  2665 => x"d0055154",
  2666 => x"80dda008",
  2667 => x"7481b72d",
  2668 => x"81195974",
  2669 => x"8b24a438",
  2670 => x"80d1d004",
  2671 => x"74902975",
  2672 => x"31701080",
  2673 => x"e4d0058c",
  2674 => x"77315751",
  2675 => x"54807481",
  2676 => x"b72d9e14",
  2677 => x"ff165654",
  2678 => x"74f33802",
  2679 => x"a4050d04",
  2680 => x"02fc050d",
  2681 => x"80dd9c08",
  2682 => x"135180d0",
  2683 => x"812d80dd",
  2684 => x"a008802e",
  2685 => x"8a3880dd",
  2686 => x"a0085180",
  2687 => x"c1812d80",
  2688 => x"0b80dd9c",
  2689 => x"0c80d18a",
  2690 => x"2daf872d",
  2691 => x"0284050d",
  2692 => x"0402fc05",
  2693 => x"0d725170",
  2694 => x"fd2eb238",
  2695 => x"70fd248b",
  2696 => x"3870fc2e",
  2697 => x"80d03880",
  2698 => x"d5800470",
  2699 => x"fe2eb938",
  2700 => x"70ff2e09",
  2701 => x"810680c8",
  2702 => x"3880dd9c",
  2703 => x"08517080",
  2704 => x"2ebe38ff",
  2705 => x"1180dd9c",
  2706 => x"0c80d580",
  2707 => x"0480dd9c",
  2708 => x"08f40570",
  2709 => x"80dd9c0c",
  2710 => x"51708025",
  2711 => x"a338800b",
  2712 => x"80dd9c0c",
  2713 => x"80d58004",
  2714 => x"80dd9c08",
  2715 => x"810580dd",
  2716 => x"9c0c80d5",
  2717 => x"800480dd",
  2718 => x"9c088c05",
  2719 => x"80dd9c0c",
  2720 => x"80d18a2d",
  2721 => x"af872d02",
  2722 => x"84050d04",
  2723 => x"02fc050d",
  2724 => x"800b80dd",
  2725 => x"9c0c80d1",
  2726 => x"8a2dae83",
  2727 => x"2d80dda0",
  2728 => x"0880dd8c",
  2729 => x"0c80dbe8",
  2730 => x"51b0ad2d",
  2731 => x"0284050d",
  2732 => x"047180e4",
  2733 => x"cc0c0400",
  2734 => x"00ffffff",
  2735 => x"ff00ffff",
  2736 => x"ffff00ff",
  2737 => x"ffffff00",
  2738 => x"30313233",
  2739 => x"34353637",
  2740 => x"38394142",
  2741 => x"43444546",
  2742 => x"00000000",
  2743 => x"52657365",
  2744 => x"74000000",
  2745 => x"5363616e",
  2746 => x"6c696e65",
  2747 => x"73000000",
  2748 => x"50414c20",
  2749 => x"2f204e54",
  2750 => x"53430000",
  2751 => x"436f6c6f",
  2752 => x"72000000",
  2753 => x"44696666",
  2754 => x"6963756c",
  2755 => x"74792041",
  2756 => x"00000000",
  2757 => x"44696666",
  2758 => x"6963756c",
  2759 => x"74792042",
  2760 => x"00000000",
  2761 => x"2a537570",
  2762 => x"65726368",
  2763 => x"69702069",
  2764 => x"6e206361",
  2765 => x"72747269",
  2766 => x"64676500",
  2767 => x"2a42616e",
  2768 => x"6b204530",
  2769 => x"00000000",
  2770 => x"2a42616e",
  2771 => x"6b204537",
  2772 => x"00000000",
  2773 => x"53656c65",
  2774 => x"63740000",
  2775 => x"53746172",
  2776 => x"74000000",
  2777 => x"4c6f6164",
  2778 => x"20524f4d",
  2779 => x"20100000",
  2780 => x"45786974",
  2781 => x"00000000",
  2782 => x"524f4d20",
  2783 => x"6c6f6164",
  2784 => x"696e6720",
  2785 => x"6661696c",
  2786 => x"65640000",
  2787 => x"4f4b0000",
  2788 => x"496e6974",
  2789 => x"69616c69",
  2790 => x"7a696e67",
  2791 => x"20534420",
  2792 => x"63617264",
  2793 => x"0a000000",
  2794 => x"16200000",
  2795 => x"14200000",
  2796 => x"15200000",
  2797 => x"53442069",
  2798 => x"6e69742e",
  2799 => x"2e2e0a00",
  2800 => x"53442063",
  2801 => x"61726420",
  2802 => x"72657365",
  2803 => x"74206661",
  2804 => x"696c6564",
  2805 => x"210a0000",
  2806 => x"53444843",
  2807 => x"20657272",
  2808 => x"6f72210a",
  2809 => x"00000000",
  2810 => x"57726974",
  2811 => x"65206661",
  2812 => x"696c6564",
  2813 => x"0a000000",
  2814 => x"52656164",
  2815 => x"20666169",
  2816 => x"6c65640a",
  2817 => x"00000000",
  2818 => x"43617264",
  2819 => x"20696e69",
  2820 => x"74206661",
  2821 => x"696c6564",
  2822 => x"0a000000",
  2823 => x"46415431",
  2824 => x"36202020",
  2825 => x"00000000",
  2826 => x"46415433",
  2827 => x"32202020",
  2828 => x"00000000",
  2829 => x"4e6f2070",
  2830 => x"61727469",
  2831 => x"74696f6e",
  2832 => x"20736967",
  2833 => x"0a000000",
  2834 => x"42616420",
  2835 => x"70617274",
  2836 => x"0a000000",
  2837 => x"4261636b",
  2838 => x"00000000",
  2839 => x"00000002",
  2840 => x"00000002",
  2841 => x"00002adc",
  2842 => x"0000035a",
  2843 => x"00000001",
  2844 => x"00002ae4",
  2845 => x"00000000",
  2846 => x"00000001",
  2847 => x"00002af0",
  2848 => x"00000001",
  2849 => x"00000001",
  2850 => x"00002afc",
  2851 => x"00000002",
  2852 => x"00000001",
  2853 => x"00002b04",
  2854 => x"00000003",
  2855 => x"00000001",
  2856 => x"00002b14",
  2857 => x"00000004",
  2858 => x"00000001",
  2859 => x"00002b24",
  2860 => x"00000005",
  2861 => x"00000001",
  2862 => x"00002b3c",
  2863 => x"00000008",
  2864 => x"00000001",
  2865 => x"00002b48",
  2866 => x"00000009",
  2867 => x"00000002",
  2868 => x"00002b54",
  2869 => x"0000036e",
  2870 => x"00000002",
  2871 => x"00002b5c",
  2872 => x"00000a3f",
  2873 => x"00000002",
  2874 => x"00002b64",
  2875 => x"00002a8c",
  2876 => x"00000002",
  2877 => x"00002b70",
  2878 => x"00001720",
  2879 => x"00000000",
  2880 => x"00000000",
  2881 => x"00000000",
  2882 => x"00000004",
  2883 => x"00002b78",
  2884 => x"00002d08",
  2885 => x"00000004",
  2886 => x"00002b8c",
  2887 => x"00002c60",
  2888 => x"00000000",
  2889 => x"00000000",
  2890 => x"00000000",
  2891 => x"00000000",
  2892 => x"00000000",
  2893 => x"00000000",
  2894 => x"00000000",
  2895 => x"00000000",
  2896 => x"00000000",
  2897 => x"00000000",
  2898 => x"00000000",
  2899 => x"00000000",
  2900 => x"00000000",
  2901 => x"00000000",
  2902 => x"00000000",
  2903 => x"00000000",
  2904 => x"00000000",
  2905 => x"00000000",
  2906 => x"00000000",
  2907 => x"761c1c1c",
  2908 => x"1c1c051c",
  2909 => x"1c1c1c1c",
  2910 => x"f2f5fafd",
  2911 => x"5a000000",
  2912 => x"00000000",
  2913 => x"00000000",
  2914 => x"00000000",
  2915 => x"00000000",
  2916 => x"00000000",
  2917 => x"00000000",
  2918 => x"00000000",
  2919 => x"00000000",
  2920 => x"00000000",
  2921 => x"00000000",
  2922 => x"00000000",
  2923 => x"00000000",
  2924 => x"00000000",
  2925 => x"00000000",
  2926 => x"00000000",
  2927 => x"00000000",
  2928 => x"00000000",
  2929 => x"00000000",
  2930 => x"0001ffff",
  2931 => x"0001ffff",
  2932 => x"0001ffff",
  2933 => x"00000000",
  2934 => x"00000000",
  2935 => x"00000006",
  2936 => x"00000000",
  2937 => x"00000000",
  2938 => x"00000002",
  2939 => x"00003250",
  2940 => x"00002850",
  2941 => x"00000002",
  2942 => x"0000326e",
  2943 => x"00002850",
  2944 => x"00000002",
  2945 => x"0000328c",
  2946 => x"00002850",
  2947 => x"00000002",
  2948 => x"000032aa",
  2949 => x"00002850",
  2950 => x"00000002",
  2951 => x"000032c8",
  2952 => x"00002850",
  2953 => x"00000002",
  2954 => x"000032e6",
  2955 => x"00002850",
  2956 => x"00000002",
  2957 => x"00003304",
  2958 => x"00002850",
  2959 => x"00000002",
  2960 => x"00003322",
  2961 => x"00002850",
  2962 => x"00000002",
  2963 => x"00003340",
  2964 => x"00002850",
  2965 => x"00000002",
  2966 => x"0000335e",
  2967 => x"00002850",
  2968 => x"00000002",
  2969 => x"0000337c",
  2970 => x"00002850",
  2971 => x"00000002",
  2972 => x"0000339a",
  2973 => x"00002850",
  2974 => x"00000002",
  2975 => x"000033b8",
  2976 => x"00002850",
  2977 => x"00000004",
  2978 => x"00002c54",
  2979 => x"00000000",
  2980 => x"00000000",
  2981 => x"00000000",
  2982 => x"00002a11",
  2983 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

