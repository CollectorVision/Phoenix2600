-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80dd",
     9 => x"a4080b0b",
    10 => x"80dda808",
    11 => x"0b0b80dd",
    12 => x"ac080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"ddac0c0b",
    16 => x"0b80dda8",
    17 => x"0c0b0b80",
    18 => x"dda40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d5bc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80dda470",
    57 => x"80e7dc27",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a6b7",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80dd",
    65 => x"b40c9f0b",
    66 => x"80ddb80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"ddb808ff",
    70 => x"0580ddb8",
    71 => x"0c80ddb8",
    72 => x"088025e8",
    73 => x"3880ddb4",
    74 => x"08ff0580",
    75 => x"ddb40c80",
    76 => x"ddb40880",
    77 => x"25d03880",
    78 => x"0b80ddb8",
    79 => x"0c800b80",
    80 => x"ddb40c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80ddb408",
   100 => x"25913882",
   101 => x"c82d80dd",
   102 => x"b408ff05",
   103 => x"80ddb40c",
   104 => x"838a0480",
   105 => x"ddb40880",
   106 => x"ddb80853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80ddb408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"ddb80881",
   116 => x"0580ddb8",
   117 => x"0c80ddb8",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80ddb8",
   121 => x"0c80ddb4",
   122 => x"08810580",
   123 => x"ddb40c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480dd",
   128 => x"b8088105",
   129 => x"80ddb80c",
   130 => x"80ddb808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80ddb8",
   134 => x"0c80ddb4",
   135 => x"08810580",
   136 => x"ddb40c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"ddbc0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"ddbc0c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280dd",
   177 => x"bc088407",
   178 => x"80ddbc0c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80d8",
   183 => x"e00c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80ddbc",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80dd",
   208 => x"a40c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02f4050d",
  1093 => x"80d8f80b",
  1094 => x"80f52d80",
  1095 => x"dbe00870",
  1096 => x"81065354",
  1097 => x"5270802e",
  1098 => x"85387184",
  1099 => x"07527281",
  1100 => x"2a708106",
  1101 => x"51517080",
  1102 => x"2e853871",
  1103 => x"82075272",
  1104 => x"822a7081",
  1105 => x"06515170",
  1106 => x"802e8538",
  1107 => x"71810752",
  1108 => x"72832a70",
  1109 => x"81065151",
  1110 => x"70802e85",
  1111 => x"38718807",
  1112 => x"5272842a",
  1113 => x"70810651",
  1114 => x"5170802e",
  1115 => x"85387190",
  1116 => x"07527285",
  1117 => x"2a708106",
  1118 => x"51517080",
  1119 => x"2e853871",
  1120 => x"a0075272",
  1121 => x"882a7081",
  1122 => x"06515170",
  1123 => x"802e8638",
  1124 => x"7180c007",
  1125 => x"5272892a",
  1126 => x"70810651",
  1127 => x"5170802e",
  1128 => x"86387181",
  1129 => x"80075271",
  1130 => x"fc0c7180",
  1131 => x"dda40c02",
  1132 => x"8c050d04",
  1133 => x"02cc050d",
  1134 => x"7e5d800b",
  1135 => x"80dbe008",
  1136 => x"81800671",
  1137 => x"5c5d5b81",
  1138 => x"0bec0c84",
  1139 => x"0bec0c7c",
  1140 => x"5280ddc0",
  1141 => x"5180cc8b",
  1142 => x"2d80dda4",
  1143 => x"087b2e80",
  1144 => x"ff3880dd",
  1145 => x"c4087bff",
  1146 => x"12575957",
  1147 => x"747b2e8b",
  1148 => x"38811875",
  1149 => x"812a5658",
  1150 => x"74f738f7",
  1151 => x"1858815b",
  1152 => x"80772580",
  1153 => x"db387752",
  1154 => x"745184a8",
  1155 => x"2d80de94",
  1156 => x"5280ddc0",
  1157 => x"5180cee0",
  1158 => x"2d80dda4",
  1159 => x"08802ea6",
  1160 => x"3880de94",
  1161 => x"597ba738",
  1162 => x"83ff5678",
  1163 => x"7081055a",
  1164 => x"80f52d7a",
  1165 => x"811c5ce4",
  1166 => x"0ce80cff",
  1167 => x"16567580",
  1168 => x"25e938a4",
  1169 => x"ce0480dd",
  1170 => x"a4085b84",
  1171 => x"805780dd",
  1172 => x"c05180ce",
  1173 => x"af2dfc80",
  1174 => x"17811656",
  1175 => x"57a48004",
  1176 => x"80ddc408",
  1177 => x"f80c881d",
  1178 => x"55807580",
  1179 => x"f52d7081",
  1180 => x"ff065558",
  1181 => x"5472742e",
  1182 => x"b6388115",
  1183 => x"80f52d53",
  1184 => x"72742eab",
  1185 => x"38738216",
  1186 => x"80f52d54",
  1187 => x"567280d3",
  1188 => x"2e098106",
  1189 => x"83388156",
  1190 => x"7280f332",
  1191 => x"70098105",
  1192 => x"70802578",
  1193 => x"07515153",
  1194 => x"72802e83",
  1195 => x"38a05480",
  1196 => x"7781ff06",
  1197 => x"54567280",
  1198 => x"c52e0981",
  1199 => x"06833881",
  1200 => x"567280e5",
  1201 => x"32700981",
  1202 => x"05708025",
  1203 => x"78075151",
  1204 => x"5372802e",
  1205 => x"a4388115",
  1206 => x"80f52d53",
  1207 => x"72b02e09",
  1208 => x"81068938",
  1209 => x"73828007",
  1210 => x"54a5f904",
  1211 => x"72b72e09",
  1212 => x"81068638",
  1213 => x"73848007",
  1214 => x"5473802e",
  1215 => x"913880db",
  1216 => x"e008f9df",
  1217 => x"06740780",
  1218 => x"dbe00ca2",
  1219 => x"902d800b",
  1220 => x"e00c8051",
  1221 => x"86da2d86",
  1222 => x"c72d7a80",
  1223 => x"2e883880",
  1224 => x"d8e451a6",
  1225 => x"aa0480da",
  1226 => x"8c51b0b2",
  1227 => x"2d7a80dd",
  1228 => x"a40c02b4",
  1229 => x"050d0402",
  1230 => x"f4050d84",
  1231 => x"0bec0c81",
  1232 => x"0be00cad",
  1233 => x"ef2da7c9",
  1234 => x"2d81f92d",
  1235 => x"8352add2",
  1236 => x"2d815185",
  1237 => x"8d2dff12",
  1238 => x"52718025",
  1239 => x"f138840b",
  1240 => x"ec0c80d7",
  1241 => x"945186a0",
  1242 => x"2d80c2b0",
  1243 => x"2d80dda4",
  1244 => x"08802ebe",
  1245 => x"38a3b451",
  1246 => x"80d5b62d",
  1247 => x"80d8e451",
  1248 => x"b0b22dae",
  1249 => x"912da8f4",
  1250 => x"2d80dda4",
  1251 => x"08810652",
  1252 => x"71802e86",
  1253 => x"38805194",
  1254 => x"bf2db0c5",
  1255 => x"2d80dda4",
  1256 => x"0852a290",
  1257 => x"2d865371",
  1258 => x"83388453",
  1259 => x"72ec0ca7",
  1260 => x"8604800b",
  1261 => x"80dda40c",
  1262 => x"028c050d",
  1263 => x"0471980c",
  1264 => x"04ffb008",
  1265 => x"80dda40c",
  1266 => x"04810bff",
  1267 => x"b00c0480",
  1268 => x"0bffb00c",
  1269 => x"0402d805",
  1270 => x"0dffb408",
  1271 => x"87ffff06",
  1272 => x"5a815480",
  1273 => x"7080dbcc",
  1274 => x"0880dbd0",
  1275 => x"0880dba8",
  1276 => x"5b59575a",
  1277 => x"58797406",
  1278 => x"75750652",
  1279 => x"5271712e",
  1280 => x"8d388077",
  1281 => x"818a2d73",
  1282 => x"09750672",
  1283 => x"07557680",
  1284 => x"e02d7083",
  1285 => x"ffff0653",
  1286 => x"517180e4",
  1287 => x"2e098106",
  1288 => x"a2387474",
  1289 => x"06707776",
  1290 => x"06327009",
  1291 => x"81057072",
  1292 => x"079f2a7b",
  1293 => x"0577097a",
  1294 => x"0674075a",
  1295 => x"5b535353",
  1296 => x"a8d10471",
  1297 => x"80e42689",
  1298 => x"38811151",
  1299 => x"7077818a",
  1300 => x"2d731081",
  1301 => x"1a821959",
  1302 => x"5a549079",
  1303 => x"25ff9638",
  1304 => x"7580dbd0",
  1305 => x"0c7480db",
  1306 => x"cc0c7780",
  1307 => x"dda40c02",
  1308 => x"a8050d04",
  1309 => x"02d0050d",
  1310 => x"805caa84",
  1311 => x"0480dda4",
  1312 => x"0881f02e",
  1313 => x"0981068a",
  1314 => x"38810b80",
  1315 => x"dbd80caa",
  1316 => x"840480dd",
  1317 => x"a40881e0",
  1318 => x"2e098106",
  1319 => x"8a38810b",
  1320 => x"80dbdc0c",
  1321 => x"aa840480",
  1322 => x"dda40852",
  1323 => x"80dbdc08",
  1324 => x"802e8938",
  1325 => x"80dda408",
  1326 => x"81800552",
  1327 => x"71842c72",
  1328 => x"8f065353",
  1329 => x"80dbd808",
  1330 => x"802e9a38",
  1331 => x"72842980",
  1332 => x"dab00572",
  1333 => x"1381712b",
  1334 => x"70097308",
  1335 => x"06730c51",
  1336 => x"5353a9f8",
  1337 => x"04728429",
  1338 => x"80dab005",
  1339 => x"72138371",
  1340 => x"2b720807",
  1341 => x"720c5353",
  1342 => x"800b80db",
  1343 => x"dc0c800b",
  1344 => x"80dbd80c",
  1345 => x"80ddcc51",
  1346 => x"acc52d80",
  1347 => x"dda408ff",
  1348 => x"24feea38",
  1349 => x"a7d52d80",
  1350 => x"dda40880",
  1351 => x"2e81b038",
  1352 => x"8159800b",
  1353 => x"80dbd408",
  1354 => x"80dbd008",
  1355 => x"80db845a",
  1356 => x"5c5c587a",
  1357 => x"79067a7a",
  1358 => x"06545271",
  1359 => x"732e80f8",
  1360 => x"38720981",
  1361 => x"05707407",
  1362 => x"802580da",
  1363 => x"f01a80f5",
  1364 => x"2d70842c",
  1365 => x"718f0658",
  1366 => x"53575752",
  1367 => x"75802ea3",
  1368 => x"38718429",
  1369 => x"80dab005",
  1370 => x"74158371",
  1371 => x"2b720807",
  1372 => x"720c5452",
  1373 => x"7680e02d",
  1374 => x"81055271",
  1375 => x"77818a2d",
  1376 => x"ab990471",
  1377 => x"842980da",
  1378 => x"b0057415",
  1379 => x"81712b70",
  1380 => x"09730806",
  1381 => x"730c5153",
  1382 => x"53748532",
  1383 => x"70098105",
  1384 => x"70802551",
  1385 => x"51527580",
  1386 => x"2e8e3881",
  1387 => x"70730653",
  1388 => x"5371802e",
  1389 => x"8338725c",
  1390 => x"78108119",
  1391 => x"82195959",
  1392 => x"59907825",
  1393 => x"feed3880",
  1394 => x"dbd00880",
  1395 => x"dbd40c7b",
  1396 => x"80dda40c",
  1397 => x"02b0050d",
  1398 => x"0402f805",
  1399 => x"0d80dab0",
  1400 => x"528f5180",
  1401 => x"72708405",
  1402 => x"540cff11",
  1403 => x"51708025",
  1404 => x"f2380288",
  1405 => x"050d0402",
  1406 => x"f0050d75",
  1407 => x"51a7cf2d",
  1408 => x"70822cfc",
  1409 => x"0680dab0",
  1410 => x"1172109e",
  1411 => x"06710870",
  1412 => x"722a7083",
  1413 => x"0682742b",
  1414 => x"70097406",
  1415 => x"760c5451",
  1416 => x"56575351",
  1417 => x"53a7c92d",
  1418 => x"7180dda4",
  1419 => x"0c029005",
  1420 => x"0d0402fc",
  1421 => x"050d7251",
  1422 => x"80710c80",
  1423 => x"0b84120c",
  1424 => x"0284050d",
  1425 => x"0402f005",
  1426 => x"0d757008",
  1427 => x"84120853",
  1428 => x"5353ff54",
  1429 => x"71712ea8",
  1430 => x"38a7cf2d",
  1431 => x"84130870",
  1432 => x"84291488",
  1433 => x"11700870",
  1434 => x"81ff0684",
  1435 => x"18088111",
  1436 => x"8706841a",
  1437 => x"0c535155",
  1438 => x"515151a7",
  1439 => x"c92d7154",
  1440 => x"7380dda4",
  1441 => x"0c029005",
  1442 => x"0d0402f8",
  1443 => x"050da7cf",
  1444 => x"2de00870",
  1445 => x"8b2a7081",
  1446 => x"06515252",
  1447 => x"70802ea1",
  1448 => x"3880ddcc",
  1449 => x"08708429",
  1450 => x"80ddd405",
  1451 => x"7381ff06",
  1452 => x"710c5151",
  1453 => x"80ddcc08",
  1454 => x"81118706",
  1455 => x"80ddcc0c",
  1456 => x"51800b80",
  1457 => x"ddf40ca7",
  1458 => x"c12da7c9",
  1459 => x"2d028805",
  1460 => x"0d0402fc",
  1461 => x"050da7cf",
  1462 => x"2d810b80",
  1463 => x"ddf40ca7",
  1464 => x"c92d80dd",
  1465 => x"f4085170",
  1466 => x"f9380284",
  1467 => x"050d0402",
  1468 => x"fc050d80",
  1469 => x"ddcc51ac",
  1470 => x"b22dabd9",
  1471 => x"2dad8a51",
  1472 => x"a7bd2d02",
  1473 => x"84050d04",
  1474 => x"80de8008",
  1475 => x"80dda40c",
  1476 => x"0402fc05",
  1477 => x"0d810b80",
  1478 => x"dbe40c81",
  1479 => x"51858d2d",
  1480 => x"0284050d",
  1481 => x"0402fc05",
  1482 => x"0daeaf04",
  1483 => x"a8f42d80",
  1484 => x"f651abf7",
  1485 => x"2d80dda4",
  1486 => x"08f23880",
  1487 => x"da51abf7",
  1488 => x"2d80dda4",
  1489 => x"08e63880",
  1490 => x"dda40880",
  1491 => x"dbe40c80",
  1492 => x"dda40851",
  1493 => x"858d2d02",
  1494 => x"84050d04",
  1495 => x"02ec050d",
  1496 => x"76548052",
  1497 => x"870b8815",
  1498 => x"80f52d56",
  1499 => x"53747224",
  1500 => x"8338a053",
  1501 => x"72518384",
  1502 => x"2d81128b",
  1503 => x"1580f52d",
  1504 => x"54527272",
  1505 => x"25de3802",
  1506 => x"94050d04",
  1507 => x"02f0050d",
  1508 => x"80de8008",
  1509 => x"5481f92d",
  1510 => x"800b80de",
  1511 => x"840c7308",
  1512 => x"802e8189",
  1513 => x"38820b80",
  1514 => x"ddb80c80",
  1515 => x"de84088f",
  1516 => x"0680ddb4",
  1517 => x"0c730852",
  1518 => x"71832e96",
  1519 => x"38718326",
  1520 => x"89387181",
  1521 => x"2eb038b0",
  1522 => x"96047185",
  1523 => x"2ea038b0",
  1524 => x"96048814",
  1525 => x"80f52d84",
  1526 => x"150880d7",
  1527 => x"ac535452",
  1528 => x"86a02d71",
  1529 => x"84291370",
  1530 => x"085252b0",
  1531 => x"9a047351",
  1532 => x"aedc2db0",
  1533 => x"960480db",
  1534 => x"e0088815",
  1535 => x"082c7081",
  1536 => x"06515271",
  1537 => x"802e8838",
  1538 => x"80d7b051",
  1539 => x"b0930480",
  1540 => x"d7b45186",
  1541 => x"a02d8414",
  1542 => x"085186a0",
  1543 => x"2d80de84",
  1544 => x"08810580",
  1545 => x"de840c8c",
  1546 => x"1454af9e",
  1547 => x"04029005",
  1548 => x"0d047180",
  1549 => x"de800caf",
  1550 => x"8c2d80de",
  1551 => x"8408ff05",
  1552 => x"80de880c",
  1553 => x"0402e805",
  1554 => x"0d80de80",
  1555 => x"0880de8c",
  1556 => x"08575580",
  1557 => x"f651abf7",
  1558 => x"2d80dda4",
  1559 => x"08812a70",
  1560 => x"81065152",
  1561 => x"71802ea4",
  1562 => x"38b0ef04",
  1563 => x"a8f42d80",
  1564 => x"f651abf7",
  1565 => x"2d80dda4",
  1566 => x"08f23880",
  1567 => x"dbe40881",
  1568 => x"327080db",
  1569 => x"e40c7052",
  1570 => x"52858d2d",
  1571 => x"800b80dd",
  1572 => x"f80c800b",
  1573 => x"80ddfc0c",
  1574 => x"80dbe408",
  1575 => x"838d3880",
  1576 => x"da51abf7",
  1577 => x"2d80dda4",
  1578 => x"08802e8c",
  1579 => x"3880ddf8",
  1580 => x"08818007",
  1581 => x"80ddf80c",
  1582 => x"80d951ab",
  1583 => x"f72d80dd",
  1584 => x"a408802e",
  1585 => x"8c3880dd",
  1586 => x"f80880c0",
  1587 => x"0780ddf8",
  1588 => x"0c819451",
  1589 => x"abf72d80",
  1590 => x"dda40880",
  1591 => x"2e8b3880",
  1592 => x"ddf80890",
  1593 => x"0780ddf8",
  1594 => x"0c819151",
  1595 => x"abf72d80",
  1596 => x"dda40880",
  1597 => x"2e8b3880",
  1598 => x"ddf808a0",
  1599 => x"0780ddf8",
  1600 => x"0c81f551",
  1601 => x"abf72d80",
  1602 => x"dda40880",
  1603 => x"2e8b3880",
  1604 => x"ddf80881",
  1605 => x"0780ddf8",
  1606 => x"0c81f251",
  1607 => x"abf72d80",
  1608 => x"dda40880",
  1609 => x"2e8b3880",
  1610 => x"ddf80882",
  1611 => x"0780ddf8",
  1612 => x"0c81eb51",
  1613 => x"abf72d80",
  1614 => x"dda40880",
  1615 => x"2e8b3880",
  1616 => x"ddf80884",
  1617 => x"0780ddf8",
  1618 => x"0c81f451",
  1619 => x"abf72d80",
  1620 => x"dda40880",
  1621 => x"2e8b3880",
  1622 => x"ddf80888",
  1623 => x"0780ddf8",
  1624 => x"0c80d851",
  1625 => x"abf72d80",
  1626 => x"dda40880",
  1627 => x"2e8c3880",
  1628 => x"ddfc0881",
  1629 => x"800780dd",
  1630 => x"fc0c9251",
  1631 => x"abf72d80",
  1632 => x"dda40880",
  1633 => x"2e8c3880",
  1634 => x"ddfc0880",
  1635 => x"c00780dd",
  1636 => x"fc0c9451",
  1637 => x"abf72d80",
  1638 => x"dda40880",
  1639 => x"2e8b3880",
  1640 => x"ddfc0890",
  1641 => x"0780ddfc",
  1642 => x"0c9151ab",
  1643 => x"f72d80dd",
  1644 => x"a408802e",
  1645 => x"8b3880dd",
  1646 => x"fc08a007",
  1647 => x"80ddfc0c",
  1648 => x"9d51abf7",
  1649 => x"2d80dda4",
  1650 => x"08802e8b",
  1651 => x"3880ddfc",
  1652 => x"08810780",
  1653 => x"ddfc0c9b",
  1654 => x"51abf72d",
  1655 => x"80dda408",
  1656 => x"802e8b38",
  1657 => x"80ddfc08",
  1658 => x"820780dd",
  1659 => x"fc0c9c51",
  1660 => x"abf72d80",
  1661 => x"dda40880",
  1662 => x"2e8b3880",
  1663 => x"ddfc0884",
  1664 => x"0780ddfc",
  1665 => x"0ca351ab",
  1666 => x"f72d80dd",
  1667 => x"a408802e",
  1668 => x"8b3880dd",
  1669 => x"fc088807",
  1670 => x"80ddfc0c",
  1671 => x"81fd51ab",
  1672 => x"f72d81fa",
  1673 => x"51abf72d",
  1674 => x"ba800481",
  1675 => x"f551abf7",
  1676 => x"2d80dda4",
  1677 => x"08812a70",
  1678 => x"81065152",
  1679 => x"71802eb3",
  1680 => x"3880de88",
  1681 => x"08527180",
  1682 => x"2e8a38ff",
  1683 => x"1280de88",
  1684 => x"0cb4f304",
  1685 => x"80de8408",
  1686 => x"1080de84",
  1687 => x"08057084",
  1688 => x"29165152",
  1689 => x"88120880",
  1690 => x"2e8938ff",
  1691 => x"51881208",
  1692 => x"52712d81",
  1693 => x"f251abf7",
  1694 => x"2d80dda4",
  1695 => x"08812a70",
  1696 => x"81065152",
  1697 => x"71802eb4",
  1698 => x"3880de84",
  1699 => x"08ff1180",
  1700 => x"de880856",
  1701 => x"53537372",
  1702 => x"258a3881",
  1703 => x"1480de88",
  1704 => x"0cb5bc04",
  1705 => x"72101370",
  1706 => x"84291651",
  1707 => x"52881208",
  1708 => x"802e8938",
  1709 => x"fe518812",
  1710 => x"0852712d",
  1711 => x"81fd51ab",
  1712 => x"f72d80dd",
  1713 => x"a408812a",
  1714 => x"70810651",
  1715 => x"5271802e",
  1716 => x"b13880de",
  1717 => x"8808802e",
  1718 => x"8a38800b",
  1719 => x"80de880c",
  1720 => x"b6820480",
  1721 => x"de840810",
  1722 => x"80de8408",
  1723 => x"05708429",
  1724 => x"16515288",
  1725 => x"1208802e",
  1726 => x"8938fd51",
  1727 => x"88120852",
  1728 => x"712d81fa",
  1729 => x"51abf72d",
  1730 => x"80dda408",
  1731 => x"812a7081",
  1732 => x"06515271",
  1733 => x"802eb138",
  1734 => x"80de8408",
  1735 => x"ff115452",
  1736 => x"80de8808",
  1737 => x"73258938",
  1738 => x"7280de88",
  1739 => x"0cb6c804",
  1740 => x"71101270",
  1741 => x"84291651",
  1742 => x"52881208",
  1743 => x"802e8938",
  1744 => x"fc518812",
  1745 => x"0852712d",
  1746 => x"80de8808",
  1747 => x"70535473",
  1748 => x"802e8a38",
  1749 => x"8c15ff15",
  1750 => x"5555b6cf",
  1751 => x"04820b80",
  1752 => x"ddb80c71",
  1753 => x"8f0680dd",
  1754 => x"b40c81eb",
  1755 => x"51abf72d",
  1756 => x"80dda408",
  1757 => x"812a7081",
  1758 => x"06515271",
  1759 => x"802ead38",
  1760 => x"7408852e",
  1761 => x"098106a4",
  1762 => x"38881580",
  1763 => x"f52dff05",
  1764 => x"52718816",
  1765 => x"81b72d71",
  1766 => x"982b5271",
  1767 => x"80258838",
  1768 => x"800b8816",
  1769 => x"81b72d74",
  1770 => x"51aedc2d",
  1771 => x"81f451ab",
  1772 => x"f72d80dd",
  1773 => x"a408812a",
  1774 => x"70810651",
  1775 => x"5271802e",
  1776 => x"b3387408",
  1777 => x"852e0981",
  1778 => x"06aa3888",
  1779 => x"1580f52d",
  1780 => x"81055271",
  1781 => x"881681b7",
  1782 => x"2d7181ff",
  1783 => x"068b1680",
  1784 => x"f52d5452",
  1785 => x"72722787",
  1786 => x"38728816",
  1787 => x"81b72d74",
  1788 => x"51aedc2d",
  1789 => x"80da51ab",
  1790 => x"f72d80dd",
  1791 => x"a408812a",
  1792 => x"70810651",
  1793 => x"5271802e",
  1794 => x"81ad3880",
  1795 => x"de800880",
  1796 => x"de880855",
  1797 => x"5373802e",
  1798 => x"8a388c13",
  1799 => x"ff155553",
  1800 => x"b8950472",
  1801 => x"08527182",
  1802 => x"2ea63871",
  1803 => x"82268938",
  1804 => x"71812eaa",
  1805 => x"38b9b704",
  1806 => x"71832eb4",
  1807 => x"3871842e",
  1808 => x"09810680",
  1809 => x"f2388813",
  1810 => x"0851b0b2",
  1811 => x"2db9b704",
  1812 => x"80de8808",
  1813 => x"51881308",
  1814 => x"52712db9",
  1815 => x"b704810b",
  1816 => x"8814082b",
  1817 => x"80dbe008",
  1818 => x"3280dbe0",
  1819 => x"0cb98b04",
  1820 => x"881380f5",
  1821 => x"2d81058b",
  1822 => x"1480f52d",
  1823 => x"53547174",
  1824 => x"24833880",
  1825 => x"54738814",
  1826 => x"81b72daf",
  1827 => x"8c2db9b7",
  1828 => x"04750880",
  1829 => x"2ea43875",
  1830 => x"0851abf7",
  1831 => x"2d80dda4",
  1832 => x"08810652",
  1833 => x"71802e8c",
  1834 => x"3880de88",
  1835 => x"08518416",
  1836 => x"0852712d",
  1837 => x"88165675",
  1838 => x"d8388054",
  1839 => x"800b80dd",
  1840 => x"b80c738f",
  1841 => x"0680ddb4",
  1842 => x"0ca05273",
  1843 => x"80de8808",
  1844 => x"2e098106",
  1845 => x"993880de",
  1846 => x"8408ff05",
  1847 => x"74327009",
  1848 => x"81057072",
  1849 => x"079f2a91",
  1850 => x"71315151",
  1851 => x"53537151",
  1852 => x"83842d81",
  1853 => x"14548e74",
  1854 => x"25c23880",
  1855 => x"dbe40852",
  1856 => x"7180dda4",
  1857 => x"0c029805",
  1858 => x"0d0402f4",
  1859 => x"050dd452",
  1860 => x"81ff720c",
  1861 => x"71085381",
  1862 => x"ff720c72",
  1863 => x"882b83fe",
  1864 => x"80067208",
  1865 => x"7081ff06",
  1866 => x"51525381",
  1867 => x"ff720c72",
  1868 => x"7107882b",
  1869 => x"72087081",
  1870 => x"ff065152",
  1871 => x"5381ff72",
  1872 => x"0c727107",
  1873 => x"882b7208",
  1874 => x"7081ff06",
  1875 => x"720780dd",
  1876 => x"a40c5253",
  1877 => x"028c050d",
  1878 => x"0402f405",
  1879 => x"0d747671",
  1880 => x"81ff06d4",
  1881 => x"0c535380",
  1882 => x"de900885",
  1883 => x"3871892b",
  1884 => x"5271982a",
  1885 => x"d40c7190",
  1886 => x"2a7081ff",
  1887 => x"06d40c51",
  1888 => x"71882a70",
  1889 => x"81ff06d4",
  1890 => x"0c517181",
  1891 => x"ff06d40c",
  1892 => x"72902a70",
  1893 => x"81ff06d4",
  1894 => x"0c51d408",
  1895 => x"7081ff06",
  1896 => x"515182b8",
  1897 => x"bf527081",
  1898 => x"ff2e0981",
  1899 => x"06943881",
  1900 => x"ff0bd40c",
  1901 => x"d4087081",
  1902 => x"ff06ff14",
  1903 => x"54515171",
  1904 => x"e5387080",
  1905 => x"dda40c02",
  1906 => x"8c050d04",
  1907 => x"02fc050d",
  1908 => x"81c75181",
  1909 => x"ff0bd40c",
  1910 => x"ff115170",
  1911 => x"8025f438",
  1912 => x"0284050d",
  1913 => x"0402f405",
  1914 => x"0d81ff0b",
  1915 => x"d40c9353",
  1916 => x"805287fc",
  1917 => x"80c151ba",
  1918 => x"d92d80dd",
  1919 => x"a4088b38",
  1920 => x"81ff0bd4",
  1921 => x"0c8153bc",
  1922 => x"9304bbcc",
  1923 => x"2dff1353",
  1924 => x"72de3872",
  1925 => x"80dda40c",
  1926 => x"028c050d",
  1927 => x"0402ec05",
  1928 => x"0d810b80",
  1929 => x"de900c84",
  1930 => x"54d00870",
  1931 => x"8f2a7081",
  1932 => x"06515153",
  1933 => x"72f33872",
  1934 => x"d00cbbcc",
  1935 => x"2d80d7b8",
  1936 => x"5186a02d",
  1937 => x"d008708f",
  1938 => x"2a708106",
  1939 => x"51515372",
  1940 => x"f338810b",
  1941 => x"d00cb153",
  1942 => x"805284d4",
  1943 => x"80c051ba",
  1944 => x"d92d80dd",
  1945 => x"a408812e",
  1946 => x"93387282",
  1947 => x"2ebf38ff",
  1948 => x"135372e4",
  1949 => x"38ff1454",
  1950 => x"73ffae38",
  1951 => x"bbcc2d83",
  1952 => x"aa52849c",
  1953 => x"80c851ba",
  1954 => x"d92d80dd",
  1955 => x"a408812e",
  1956 => x"09810693",
  1957 => x"38ba8a2d",
  1958 => x"80dda408",
  1959 => x"83ffff06",
  1960 => x"537283aa",
  1961 => x"2e9f38bb",
  1962 => x"e52dbdc0",
  1963 => x"0480d7c4",
  1964 => x"5186a02d",
  1965 => x"8053bf95",
  1966 => x"0480d7dc",
  1967 => x"5186a02d",
  1968 => x"8054bee6",
  1969 => x"0481ff0b",
  1970 => x"d40cb154",
  1971 => x"bbcc2d8f",
  1972 => x"cf538052",
  1973 => x"87fc80f7",
  1974 => x"51bad92d",
  1975 => x"80dda408",
  1976 => x"5580dda4",
  1977 => x"08812e09",
  1978 => x"81069c38",
  1979 => x"81ff0bd4",
  1980 => x"0c820a52",
  1981 => x"849c80e9",
  1982 => x"51bad92d",
  1983 => x"80dda408",
  1984 => x"802e8d38",
  1985 => x"bbcc2dff",
  1986 => x"135372c6",
  1987 => x"38bed904",
  1988 => x"81ff0bd4",
  1989 => x"0c80dda4",
  1990 => x"085287fc",
  1991 => x"80fa51ba",
  1992 => x"d92d80dd",
  1993 => x"a408b238",
  1994 => x"81ff0bd4",
  1995 => x"0cd40853",
  1996 => x"81ff0bd4",
  1997 => x"0c81ff0b",
  1998 => x"d40c81ff",
  1999 => x"0bd40c81",
  2000 => x"ff0bd40c",
  2001 => x"72862a70",
  2002 => x"81067656",
  2003 => x"51537296",
  2004 => x"3880dda4",
  2005 => x"0854bee6",
  2006 => x"0473822e",
  2007 => x"fedb38ff",
  2008 => x"145473fe",
  2009 => x"e7387380",
  2010 => x"de900c73",
  2011 => x"8b388152",
  2012 => x"87fc80d0",
  2013 => x"51bad92d",
  2014 => x"81ff0bd4",
  2015 => x"0cd00870",
  2016 => x"8f2a7081",
  2017 => x"06515153",
  2018 => x"72f33872",
  2019 => x"d00c81ff",
  2020 => x"0bd40c81",
  2021 => x"537280dd",
  2022 => x"a40c0294",
  2023 => x"050d0402",
  2024 => x"e8050d78",
  2025 => x"55805681",
  2026 => x"ff0bd40c",
  2027 => x"d008708f",
  2028 => x"2a708106",
  2029 => x"51515372",
  2030 => x"f3388281",
  2031 => x"0bd00c81",
  2032 => x"ff0bd40c",
  2033 => x"775287fc",
  2034 => x"80d151ba",
  2035 => x"d92d80db",
  2036 => x"c6df5480",
  2037 => x"dda40880",
  2038 => x"2e8c3880",
  2039 => x"d7fc5186",
  2040 => x"a02d80c0",
  2041 => x"bb0481ff",
  2042 => x"0bd40cd4",
  2043 => x"087081ff",
  2044 => x"06515372",
  2045 => x"81fe2e09",
  2046 => x"81069f38",
  2047 => x"80ff53ba",
  2048 => x"8a2d80dd",
  2049 => x"a4087570",
  2050 => x"8405570c",
  2051 => x"ff135372",
  2052 => x"8025ec38",
  2053 => x"815680c0",
  2054 => x"a004ff14",
  2055 => x"5473c738",
  2056 => x"81ff0bd4",
  2057 => x"0c81ff0b",
  2058 => x"d40cd008",
  2059 => x"708f2a70",
  2060 => x"81065151",
  2061 => x"5372f338",
  2062 => x"72d00c75",
  2063 => x"80dda40c",
  2064 => x"0298050d",
  2065 => x"0402e805",
  2066 => x"0d77797b",
  2067 => x"58555580",
  2068 => x"53727625",
  2069 => x"a5387470",
  2070 => x"81055680",
  2071 => x"f52d7470",
  2072 => x"81055680",
  2073 => x"f52d5252",
  2074 => x"71712e87",
  2075 => x"38815180",
  2076 => x"c0fc0481",
  2077 => x"135380c0",
  2078 => x"d1048051",
  2079 => x"7080dda4",
  2080 => x"0c029805",
  2081 => x"0d0402ec",
  2082 => x"050d7655",
  2083 => x"74802e80",
  2084 => x"c4389a15",
  2085 => x"80e02d51",
  2086 => x"80cfba2d",
  2087 => x"80dda408",
  2088 => x"80dda408",
  2089 => x"80e4c40c",
  2090 => x"80dda408",
  2091 => x"545480e4",
  2092 => x"a008802e",
  2093 => x"9b389415",
  2094 => x"80e02d51",
  2095 => x"80cfba2d",
  2096 => x"80dda408",
  2097 => x"902b83ff",
  2098 => x"f00a0670",
  2099 => x"75075153",
  2100 => x"7280e4c4",
  2101 => x"0c80e4c4",
  2102 => x"08537280",
  2103 => x"2e9e3880",
  2104 => x"e49808fe",
  2105 => x"14712980",
  2106 => x"e4ac0805",
  2107 => x"80e4c80c",
  2108 => x"70842b80",
  2109 => x"e4a40c54",
  2110 => x"80c2ab04",
  2111 => x"80e4b008",
  2112 => x"80e4c40c",
  2113 => x"80e4b408",
  2114 => x"80e4c80c",
  2115 => x"80e4a008",
  2116 => x"802e8c38",
  2117 => x"80e49808",
  2118 => x"842b5380",
  2119 => x"c2a60480",
  2120 => x"e4b80884",
  2121 => x"2b537280",
  2122 => x"e4a40c02",
  2123 => x"94050d04",
  2124 => x"02d8050d",
  2125 => x"800b80e4",
  2126 => x"a00c8454",
  2127 => x"bc9d2d80",
  2128 => x"dda40880",
  2129 => x"2e983880",
  2130 => x"de945280",
  2131 => x"51bf9f2d",
  2132 => x"80dda408",
  2133 => x"802e8738",
  2134 => x"fe5480c2",
  2135 => x"e604ff14",
  2136 => x"54738024",
  2137 => x"d738738e",
  2138 => x"3880d88c",
  2139 => x"5186a02d",
  2140 => x"735580c8",
  2141 => x"c9048056",
  2142 => x"810b80e4",
  2143 => x"cc0c8853",
  2144 => x"80d8a052",
  2145 => x"80deca51",
  2146 => x"80c0c52d",
  2147 => x"80dda408",
  2148 => x"762e0981",
  2149 => x"06893880",
  2150 => x"dda40880",
  2151 => x"e4cc0c88",
  2152 => x"5380d8ac",
  2153 => x"5280dee6",
  2154 => x"5180c0c5",
  2155 => x"2d80dda4",
  2156 => x"08893880",
  2157 => x"dda40880",
  2158 => x"e4cc0c80",
  2159 => x"e4cc0880",
  2160 => x"2e818438",
  2161 => x"80e1da0b",
  2162 => x"80f52d80",
  2163 => x"e1db0b80",
  2164 => x"f52d7198",
  2165 => x"2b71902b",
  2166 => x"0780e1dc",
  2167 => x"0b80f52d",
  2168 => x"70882b72",
  2169 => x"0780e1dd",
  2170 => x"0b80f52d",
  2171 => x"710780e2",
  2172 => x"920b80f5",
  2173 => x"2d80e293",
  2174 => x"0b80f52d",
  2175 => x"71882b07",
  2176 => x"535f5452",
  2177 => x"5a565755",
  2178 => x"7381abaa",
  2179 => x"2e098106",
  2180 => x"90387551",
  2181 => x"80cf892d",
  2182 => x"80dda408",
  2183 => x"5680c4b0",
  2184 => x"047382d4",
  2185 => x"d52e8938",
  2186 => x"80d8b851",
  2187 => x"80c4ff04",
  2188 => x"80de9452",
  2189 => x"7551bf9f",
  2190 => x"2d80dda4",
  2191 => x"085580dd",
  2192 => x"a408802e",
  2193 => x"84833888",
  2194 => x"5380d8ac",
  2195 => x"5280dee6",
  2196 => x"5180c0c5",
  2197 => x"2d80dda4",
  2198 => x"088b3881",
  2199 => x"0b80e4a0",
  2200 => x"0c80c586",
  2201 => x"04885380",
  2202 => x"d8a05280",
  2203 => x"deca5180",
  2204 => x"c0c52d80",
  2205 => x"dda40880",
  2206 => x"2e8c3880",
  2207 => x"d8cc5186",
  2208 => x"a02d80c5",
  2209 => x"e50480e2",
  2210 => x"920b80f5",
  2211 => x"2d547380",
  2212 => x"d52e0981",
  2213 => x"0680ce38",
  2214 => x"80e2930b",
  2215 => x"80f52d54",
  2216 => x"7381aa2e",
  2217 => x"098106bd",
  2218 => x"38800b80",
  2219 => x"de940b80",
  2220 => x"f52d5654",
  2221 => x"7481e92e",
  2222 => x"83388154",
  2223 => x"7481eb2e",
  2224 => x"8c388055",
  2225 => x"73752e09",
  2226 => x"810682fd",
  2227 => x"3880de9f",
  2228 => x"0b80f52d",
  2229 => x"55748e38",
  2230 => x"80dea00b",
  2231 => x"80f52d54",
  2232 => x"73822e87",
  2233 => x"38805580",
  2234 => x"c8c90480",
  2235 => x"dea10b80",
  2236 => x"f52d7080",
  2237 => x"e4980cff",
  2238 => x"0580e49c",
  2239 => x"0c80dea2",
  2240 => x"0b80f52d",
  2241 => x"80dea30b",
  2242 => x"80f52d58",
  2243 => x"76057782",
  2244 => x"80290570",
  2245 => x"80e4a80c",
  2246 => x"80dea40b",
  2247 => x"80f52d70",
  2248 => x"80e4bc0c",
  2249 => x"80e4a008",
  2250 => x"59575876",
  2251 => x"802e81b9",
  2252 => x"38885380",
  2253 => x"d8ac5280",
  2254 => x"dee65180",
  2255 => x"c0c52d80",
  2256 => x"dda40882",
  2257 => x"843880e4",
  2258 => x"98087084",
  2259 => x"2b80e4a4",
  2260 => x"0c7080e4",
  2261 => x"b80c80de",
  2262 => x"b90b80f5",
  2263 => x"2d80deb8",
  2264 => x"0b80f52d",
  2265 => x"71828029",
  2266 => x"0580deba",
  2267 => x"0b80f52d",
  2268 => x"70848080",
  2269 => x"291280de",
  2270 => x"bb0b80f5",
  2271 => x"2d708180",
  2272 => x"0a291270",
  2273 => x"80e4c00c",
  2274 => x"80e4bc08",
  2275 => x"712980e4",
  2276 => x"a8080570",
  2277 => x"80e4ac0c",
  2278 => x"80dec10b",
  2279 => x"80f52d80",
  2280 => x"dec00b80",
  2281 => x"f52d7182",
  2282 => x"80290580",
  2283 => x"dec20b80",
  2284 => x"f52d7084",
  2285 => x"80802912",
  2286 => x"80dec30b",
  2287 => x"80f52d70",
  2288 => x"982b81f0",
  2289 => x"0a067205",
  2290 => x"7080e4b0",
  2291 => x"0cfe117e",
  2292 => x"29770580",
  2293 => x"e4b40c52",
  2294 => x"59524354",
  2295 => x"5e515259",
  2296 => x"525d5759",
  2297 => x"5780c8c1",
  2298 => x"0480dea6",
  2299 => x"0b80f52d",
  2300 => x"80dea50b",
  2301 => x"80f52d71",
  2302 => x"82802905",
  2303 => x"7080e4a4",
  2304 => x"0c70a029",
  2305 => x"83ff0570",
  2306 => x"892a7080",
  2307 => x"e4b80c80",
  2308 => x"deab0b80",
  2309 => x"f52d80de",
  2310 => x"aa0b80f5",
  2311 => x"2d718280",
  2312 => x"29057080",
  2313 => x"e4c00c7b",
  2314 => x"71291e70",
  2315 => x"80e4b40c",
  2316 => x"7d80e4b0",
  2317 => x"0c730580",
  2318 => x"e4ac0c55",
  2319 => x"5e515155",
  2320 => x"55805180",
  2321 => x"c1862d81",
  2322 => x"557480dd",
  2323 => x"a40c02a8",
  2324 => x"050d0402",
  2325 => x"ec050d76",
  2326 => x"70872c71",
  2327 => x"80ff0655",
  2328 => x"565480e4",
  2329 => x"a0088a38",
  2330 => x"73882c74",
  2331 => x"81ff0654",
  2332 => x"5580de94",
  2333 => x"5280e4a8",
  2334 => x"081551bf",
  2335 => x"9f2d80dd",
  2336 => x"a4085480",
  2337 => x"dda40880",
  2338 => x"2ebb3880",
  2339 => x"e4a00880",
  2340 => x"2e9c3872",
  2341 => x"842980de",
  2342 => x"94057008",
  2343 => x"525380cf",
  2344 => x"892d80dd",
  2345 => x"a408f00a",
  2346 => x"065380c9",
  2347 => x"c3047210",
  2348 => x"80de9405",
  2349 => x"7080e02d",
  2350 => x"525380cf",
  2351 => x"ba2d80dd",
  2352 => x"a4085372",
  2353 => x"547380dd",
  2354 => x"a40c0294",
  2355 => x"050d0402",
  2356 => x"e0050d79",
  2357 => x"70842c80",
  2358 => x"e4c80805",
  2359 => x"718f0652",
  2360 => x"5553728a",
  2361 => x"3880de94",
  2362 => x"527351bf",
  2363 => x"9f2d72a0",
  2364 => x"2980de94",
  2365 => x"05548074",
  2366 => x"80f52d56",
  2367 => x"5374732e",
  2368 => x"83388153",
  2369 => x"7481e52e",
  2370 => x"81f53881",
  2371 => x"70740654",
  2372 => x"5872802e",
  2373 => x"81e9388b",
  2374 => x"1480f52d",
  2375 => x"70832a79",
  2376 => x"06585676",
  2377 => x"9c3880db",
  2378 => x"e8085372",
  2379 => x"89387280",
  2380 => x"e2940b81",
  2381 => x"b72d7680",
  2382 => x"dbe80c73",
  2383 => x"5380cc81",
  2384 => x"04758f2e",
  2385 => x"09810681",
  2386 => x"b638749f",
  2387 => x"068d2980",
  2388 => x"e2871151",
  2389 => x"53811480",
  2390 => x"f52d7370",
  2391 => x"81055581",
  2392 => x"b72d8314",
  2393 => x"80f52d73",
  2394 => x"70810555",
  2395 => x"81b72d85",
  2396 => x"1480f52d",
  2397 => x"73708105",
  2398 => x"5581b72d",
  2399 => x"871480f5",
  2400 => x"2d737081",
  2401 => x"055581b7",
  2402 => x"2d891480",
  2403 => x"f52d7370",
  2404 => x"81055581",
  2405 => x"b72d8e14",
  2406 => x"80f52d73",
  2407 => x"70810555",
  2408 => x"81b72d90",
  2409 => x"1480f52d",
  2410 => x"73708105",
  2411 => x"5581b72d",
  2412 => x"921480f5",
  2413 => x"2d737081",
  2414 => x"055581b7",
  2415 => x"2d941480",
  2416 => x"f52d7370",
  2417 => x"81055581",
  2418 => x"b72d9614",
  2419 => x"80f52d73",
  2420 => x"70810555",
  2421 => x"81b72d98",
  2422 => x"1480f52d",
  2423 => x"73708105",
  2424 => x"5581b72d",
  2425 => x"9c1480f5",
  2426 => x"2d737081",
  2427 => x"055581b7",
  2428 => x"2d9e1480",
  2429 => x"f52d7381",
  2430 => x"b72d7780",
  2431 => x"dbe80c80",
  2432 => x"537280dd",
  2433 => x"a40c02a0",
  2434 => x"050d0402",
  2435 => x"cc050d7e",
  2436 => x"605e5a80",
  2437 => x"0b80e4c4",
  2438 => x"0880e4c8",
  2439 => x"08595c56",
  2440 => x"805880e4",
  2441 => x"a408782e",
  2442 => x"81bd3877",
  2443 => x"8f06a017",
  2444 => x"57547391",
  2445 => x"3880de94",
  2446 => x"52765181",
  2447 => x"1757bf9f",
  2448 => x"2d80de94",
  2449 => x"56807680",
  2450 => x"f52d5654",
  2451 => x"74742e83",
  2452 => x"38815474",
  2453 => x"81e52e81",
  2454 => x"82388170",
  2455 => x"7506555c",
  2456 => x"73802e80",
  2457 => x"f6388b16",
  2458 => x"80f52d98",
  2459 => x"06597880",
  2460 => x"ea388b53",
  2461 => x"7c527551",
  2462 => x"80c0c52d",
  2463 => x"80dda408",
  2464 => x"80d9389c",
  2465 => x"16085180",
  2466 => x"cf892d80",
  2467 => x"dda40884",
  2468 => x"1b0c9a16",
  2469 => x"80e02d51",
  2470 => x"80cfba2d",
  2471 => x"80dda408",
  2472 => x"80dda408",
  2473 => x"881c0c80",
  2474 => x"dda40855",
  2475 => x"5580e4a0",
  2476 => x"08802e9a",
  2477 => x"38941680",
  2478 => x"e02d5180",
  2479 => x"cfba2d80",
  2480 => x"dda40890",
  2481 => x"2b83fff0",
  2482 => x"0a067016",
  2483 => x"51547388",
  2484 => x"1b0c787a",
  2485 => x"0c7b5480",
  2486 => x"cea50481",
  2487 => x"185880e4",
  2488 => x"a4087826",
  2489 => x"fec53880",
  2490 => x"e4a00880",
  2491 => x"2eb5387a",
  2492 => x"5180c8d3",
  2493 => x"2d80dda4",
  2494 => x"0880dda4",
  2495 => x"0880ffff",
  2496 => x"fff80655",
  2497 => x"5b7380ff",
  2498 => x"fffff82e",
  2499 => x"963880dd",
  2500 => x"a408fe05",
  2501 => x"80e49808",
  2502 => x"2980e4ac",
  2503 => x"08055780",
  2504 => x"cca00480",
  2505 => x"547380dd",
  2506 => x"a40c02b4",
  2507 => x"050d0402",
  2508 => x"f4050d74",
  2509 => x"70088105",
  2510 => x"710c7008",
  2511 => x"80e49c08",
  2512 => x"06535371",
  2513 => x"90388813",
  2514 => x"085180c8",
  2515 => x"d32d80dd",
  2516 => x"a4088814",
  2517 => x"0c810b80",
  2518 => x"dda40c02",
  2519 => x"8c050d04",
  2520 => x"02f0050d",
  2521 => x"75881108",
  2522 => x"fe0580e4",
  2523 => x"98082980",
  2524 => x"e4ac0811",
  2525 => x"720880e4",
  2526 => x"9c080605",
  2527 => x"79555354",
  2528 => x"54bf9f2d",
  2529 => x"0290050d",
  2530 => x"0402f405",
  2531 => x"0d747088",
  2532 => x"2a83fe80",
  2533 => x"06707298",
  2534 => x"2a077288",
  2535 => x"2b87fc80",
  2536 => x"80067398",
  2537 => x"2b81f00a",
  2538 => x"06717307",
  2539 => x"0780dda4",
  2540 => x"0c565153",
  2541 => x"51028c05",
  2542 => x"0d0402f8",
  2543 => x"050d028e",
  2544 => x"0580f52d",
  2545 => x"74882b07",
  2546 => x"7083ffff",
  2547 => x"0680dda4",
  2548 => x"0c510288",
  2549 => x"050d0402",
  2550 => x"f4050d74",
  2551 => x"76785354",
  2552 => x"52807125",
  2553 => x"97387270",
  2554 => x"81055480",
  2555 => x"f52d7270",
  2556 => x"81055481",
  2557 => x"b72dff11",
  2558 => x"5170eb38",
  2559 => x"807281b7",
  2560 => x"2d028c05",
  2561 => x"0d0402e8",
  2562 => x"050d7756",
  2563 => x"80705654",
  2564 => x"737624b7",
  2565 => x"3880e4a4",
  2566 => x"08742eaf",
  2567 => x"38735180",
  2568 => x"c9cf2d80",
  2569 => x"dda40880",
  2570 => x"dda40809",
  2571 => x"81057080",
  2572 => x"dda40807",
  2573 => x"9f2a7705",
  2574 => x"81175757",
  2575 => x"53537476",
  2576 => x"24893880",
  2577 => x"e4a40874",
  2578 => x"26d33872",
  2579 => x"80dda40c",
  2580 => x"0298050d",
  2581 => x"0402f005",
  2582 => x"0d80dda0",
  2583 => x"08165180",
  2584 => x"d0862d80",
  2585 => x"dda40880",
  2586 => x"2ea0388b",
  2587 => x"5380dda4",
  2588 => x"085280e2",
  2589 => x"945180cf",
  2590 => x"d72d80e4",
  2591 => x"d0085473",
  2592 => x"802e8738",
  2593 => x"80e29451",
  2594 => x"732d0290",
  2595 => x"050d0402",
  2596 => x"dc050d80",
  2597 => x"705a5574",
  2598 => x"80dda008",
  2599 => x"25b53880",
  2600 => x"e4a40875",
  2601 => x"2ead3878",
  2602 => x"5180c9cf",
  2603 => x"2d80dda4",
  2604 => x"08098105",
  2605 => x"7080dda4",
  2606 => x"08079f2a",
  2607 => x"7605811b",
  2608 => x"5b565474",
  2609 => x"80dda008",
  2610 => x"25893880",
  2611 => x"e4a40879",
  2612 => x"26d53880",
  2613 => x"557880e4",
  2614 => x"a4082781",
  2615 => x"e4387851",
  2616 => x"80c9cf2d",
  2617 => x"80dda408",
  2618 => x"802e81b4",
  2619 => x"3880dda4",
  2620 => x"088b0580",
  2621 => x"f52d7084",
  2622 => x"2a708106",
  2623 => x"77107884",
  2624 => x"2b80e294",
  2625 => x"0b80f52d",
  2626 => x"5c5c5351",
  2627 => x"55567380",
  2628 => x"2e80ce38",
  2629 => x"7416822b",
  2630 => x"80d3e50b",
  2631 => x"80dbf412",
  2632 => x"0c547775",
  2633 => x"311080e4",
  2634 => x"d4115556",
  2635 => x"90747081",
  2636 => x"055681b7",
  2637 => x"2da07481",
  2638 => x"b72d7681",
  2639 => x"ff068116",
  2640 => x"58547380",
  2641 => x"2e8b389c",
  2642 => x"5380e294",
  2643 => x"5280d2d8",
  2644 => x"048b5380",
  2645 => x"dda40852",
  2646 => x"80e4d616",
  2647 => x"5180d396",
  2648 => x"04741682",
  2649 => x"2b80d0d5",
  2650 => x"0b80dbf4",
  2651 => x"120c5476",
  2652 => x"81ff0681",
  2653 => x"16585473",
  2654 => x"802e8b38",
  2655 => x"9c5380e2",
  2656 => x"945280d3",
  2657 => x"8d048b53",
  2658 => x"80dda408",
  2659 => x"52777531",
  2660 => x"1080e4d4",
  2661 => x"05517655",
  2662 => x"80cfd72d",
  2663 => x"80d3b504",
  2664 => x"74902975",
  2665 => x"31701080",
  2666 => x"e4d40551",
  2667 => x"5480dda4",
  2668 => x"087481b7",
  2669 => x"2d811959",
  2670 => x"748b24a4",
  2671 => x"3880d1d5",
  2672 => x"04749029",
  2673 => x"75317010",
  2674 => x"80e4d405",
  2675 => x"8c773157",
  2676 => x"51548074",
  2677 => x"81b72d9e",
  2678 => x"14ff1656",
  2679 => x"5474f338",
  2680 => x"02a4050d",
  2681 => x"0402fc05",
  2682 => x"0d80dda0",
  2683 => x"08135180",
  2684 => x"d0862d80",
  2685 => x"dda40880",
  2686 => x"2e8a3880",
  2687 => x"dda40851",
  2688 => x"80c1862d",
  2689 => x"800b80dd",
  2690 => x"a00c80d1",
  2691 => x"8f2daf8c",
  2692 => x"2d028405",
  2693 => x"0d0402fc",
  2694 => x"050d7251",
  2695 => x"70fd2eb2",
  2696 => x"3870fd24",
  2697 => x"8b3870fc",
  2698 => x"2e80d038",
  2699 => x"80d58504",
  2700 => x"70fe2eb9",
  2701 => x"3870ff2e",
  2702 => x"09810680",
  2703 => x"c83880dd",
  2704 => x"a0085170",
  2705 => x"802ebe38",
  2706 => x"ff1180dd",
  2707 => x"a00c80d5",
  2708 => x"850480dd",
  2709 => x"a008f405",
  2710 => x"7080dda0",
  2711 => x"0c517080",
  2712 => x"25a33880",
  2713 => x"0b80dda0",
  2714 => x"0c80d585",
  2715 => x"0480dda0",
  2716 => x"08810580",
  2717 => x"dda00c80",
  2718 => x"d5850480",
  2719 => x"dda0088c",
  2720 => x"0580dda0",
  2721 => x"0c80d18f",
  2722 => x"2daf8c2d",
  2723 => x"0284050d",
  2724 => x"0402fc05",
  2725 => x"0d800b80",
  2726 => x"dda00c80",
  2727 => x"d18f2dae",
  2728 => x"882d80dd",
  2729 => x"a40880dd",
  2730 => x"900c80db",
  2731 => x"ec51b0b2",
  2732 => x"2d028405",
  2733 => x"0d047180",
  2734 => x"e4d00c04",
  2735 => x"00ffffff",
  2736 => x"ff00ffff",
  2737 => x"ffff00ff",
  2738 => x"ffffff00",
  2739 => x"30313233",
  2740 => x"34353637",
  2741 => x"38394142",
  2742 => x"43444546",
  2743 => x"00000000",
  2744 => x"52657365",
  2745 => x"74000000",
  2746 => x"5363616e",
  2747 => x"6c696e65",
  2748 => x"73000000",
  2749 => x"50414c20",
  2750 => x"2f204e54",
  2751 => x"53430000",
  2752 => x"436f6c6f",
  2753 => x"72000000",
  2754 => x"44696666",
  2755 => x"6963756c",
  2756 => x"74792041",
  2757 => x"00000000",
  2758 => x"44696666",
  2759 => x"6963756c",
  2760 => x"74792042",
  2761 => x"00000000",
  2762 => x"2a537570",
  2763 => x"65726368",
  2764 => x"69702069",
  2765 => x"6e206361",
  2766 => x"72747269",
  2767 => x"64676500",
  2768 => x"2a42616e",
  2769 => x"6b204530",
  2770 => x"00000000",
  2771 => x"2a42616e",
  2772 => x"6b204537",
  2773 => x"00000000",
  2774 => x"53656c65",
  2775 => x"63740000",
  2776 => x"53746172",
  2777 => x"74000000",
  2778 => x"4c6f6164",
  2779 => x"20524f4d",
  2780 => x"20100000",
  2781 => x"45786974",
  2782 => x"00000000",
  2783 => x"524f4d20",
  2784 => x"6c6f6164",
  2785 => x"696e6720",
  2786 => x"6661696c",
  2787 => x"65640000",
  2788 => x"4f4b0000",
  2789 => x"496e6974",
  2790 => x"69616c69",
  2791 => x"7a696e67",
  2792 => x"20534420",
  2793 => x"63617264",
  2794 => x"0a000000",
  2795 => x"16200000",
  2796 => x"14200000",
  2797 => x"15200000",
  2798 => x"53442069",
  2799 => x"6e69742e",
  2800 => x"2e2e0a00",
  2801 => x"53442063",
  2802 => x"61726420",
  2803 => x"72657365",
  2804 => x"74206661",
  2805 => x"696c6564",
  2806 => x"210a0000",
  2807 => x"53444843",
  2808 => x"20657272",
  2809 => x"6f72210a",
  2810 => x"00000000",
  2811 => x"57726974",
  2812 => x"65206661",
  2813 => x"696c6564",
  2814 => x"0a000000",
  2815 => x"52656164",
  2816 => x"20666169",
  2817 => x"6c65640a",
  2818 => x"00000000",
  2819 => x"43617264",
  2820 => x"20696e69",
  2821 => x"74206661",
  2822 => x"696c6564",
  2823 => x"0a000000",
  2824 => x"46415431",
  2825 => x"36202020",
  2826 => x"00000000",
  2827 => x"46415433",
  2828 => x"32202020",
  2829 => x"00000000",
  2830 => x"4e6f2070",
  2831 => x"61727469",
  2832 => x"74696f6e",
  2833 => x"20736967",
  2834 => x"0a000000",
  2835 => x"42616420",
  2836 => x"70617274",
  2837 => x"0a000000",
  2838 => x"4261636b",
  2839 => x"00000000",
  2840 => x"00000002",
  2841 => x"00000002",
  2842 => x"00002ae0",
  2843 => x"0000035a",
  2844 => x"00000001",
  2845 => x"00002ae8",
  2846 => x"00000000",
  2847 => x"00000001",
  2848 => x"00002af4",
  2849 => x"00000001",
  2850 => x"00000001",
  2851 => x"00002b00",
  2852 => x"00000002",
  2853 => x"00000001",
  2854 => x"00002b08",
  2855 => x"00000003",
  2856 => x"00000001",
  2857 => x"00002b18",
  2858 => x"00000004",
  2859 => x"00000001",
  2860 => x"00002b28",
  2861 => x"00000005",
  2862 => x"00000001",
  2863 => x"00002b40",
  2864 => x"00000008",
  2865 => x"00000001",
  2866 => x"00002b4c",
  2867 => x"00000009",
  2868 => x"00000002",
  2869 => x"00002b58",
  2870 => x"0000036e",
  2871 => x"00000002",
  2872 => x"00002b60",
  2873 => x"00000a3f",
  2874 => x"00000002",
  2875 => x"00002b68",
  2876 => x"00002a91",
  2877 => x"00000002",
  2878 => x"00002b74",
  2879 => x"00001725",
  2880 => x"00000000",
  2881 => x"00000000",
  2882 => x"00000000",
  2883 => x"00000004",
  2884 => x"00002b7c",
  2885 => x"00002d0c",
  2886 => x"00000004",
  2887 => x"00002b90",
  2888 => x"00002c64",
  2889 => x"00000000",
  2890 => x"00000000",
  2891 => x"00000000",
  2892 => x"00000000",
  2893 => x"00000000",
  2894 => x"00000000",
  2895 => x"00000000",
  2896 => x"00000000",
  2897 => x"00000000",
  2898 => x"00000000",
  2899 => x"00000000",
  2900 => x"00000000",
  2901 => x"00000000",
  2902 => x"00000000",
  2903 => x"00000000",
  2904 => x"00000000",
  2905 => x"00000000",
  2906 => x"00000000",
  2907 => x"00000000",
  2908 => x"761c1c1c",
  2909 => x"1c1c051c",
  2910 => x"1c1c1c1c",
  2911 => x"f2f5fafd",
  2912 => x"5a000000",
  2913 => x"00000000",
  2914 => x"00000000",
  2915 => x"00000000",
  2916 => x"00000000",
  2917 => x"00000000",
  2918 => x"00000000",
  2919 => x"00000000",
  2920 => x"00000000",
  2921 => x"00000000",
  2922 => x"00000000",
  2923 => x"00000000",
  2924 => x"00000000",
  2925 => x"00000000",
  2926 => x"00000000",
  2927 => x"00000000",
  2928 => x"00000000",
  2929 => x"00000000",
  2930 => x"00000000",
  2931 => x"0001ffff",
  2932 => x"0001ffff",
  2933 => x"0001ffff",
  2934 => x"00000000",
  2935 => x"00000000",
  2936 => x"00000006",
  2937 => x"00000000",
  2938 => x"00000000",
  2939 => x"00000002",
  2940 => x"00003254",
  2941 => x"00002855",
  2942 => x"00000002",
  2943 => x"00003272",
  2944 => x"00002855",
  2945 => x"00000002",
  2946 => x"00003290",
  2947 => x"00002855",
  2948 => x"00000002",
  2949 => x"000032ae",
  2950 => x"00002855",
  2951 => x"00000002",
  2952 => x"000032cc",
  2953 => x"00002855",
  2954 => x"00000002",
  2955 => x"000032ea",
  2956 => x"00002855",
  2957 => x"00000002",
  2958 => x"00003308",
  2959 => x"00002855",
  2960 => x"00000002",
  2961 => x"00003326",
  2962 => x"00002855",
  2963 => x"00000002",
  2964 => x"00003344",
  2965 => x"00002855",
  2966 => x"00000002",
  2967 => x"00003362",
  2968 => x"00002855",
  2969 => x"00000002",
  2970 => x"00003380",
  2971 => x"00002855",
  2972 => x"00000002",
  2973 => x"0000339e",
  2974 => x"00002855",
  2975 => x"00000002",
  2976 => x"000033bc",
  2977 => x"00002855",
  2978 => x"00000004",
  2979 => x"00002c58",
  2980 => x"00000000",
  2981 => x"00000000",
  2982 => x"00000000",
  2983 => x"00002a16",
  2984 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

