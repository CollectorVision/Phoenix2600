-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80db",
     9 => x"f0080b0b",
    10 => x"80dbf408",
    11 => x"0b0b80db",
    12 => x"f8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"dbf80c0b",
    16 => x"0b80dbf4",
    17 => x"0c0b0b80",
    18 => x"dbf00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d4c4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80dbf070",
    57 => x"80e7b027",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a7ce",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80dc",
    65 => x"800c9f0b",
    66 => x"80dc840c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"dc8408ff",
    70 => x"0580dc84",
    71 => x"0c80dc84",
    72 => x"088025e8",
    73 => x"3880dc80",
    74 => x"08ff0580",
    75 => x"dc800c80",
    76 => x"dc800880",
    77 => x"25d03880",
    78 => x"0b80dc84",
    79 => x"0c800b80",
    80 => x"dc800c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80dc8008",
   100 => x"25913882",
   101 => x"c82d80dc",
   102 => x"8008ff05",
   103 => x"80dc800c",
   104 => x"838a0480",
   105 => x"dc800880",
   106 => x"dc840853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80dc8008",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"dc840881",
   116 => x"0580dc84",
   117 => x"0c80dc84",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80dc84",
   121 => x"0c80dc80",
   122 => x"08810580",
   123 => x"dc800c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480dc",
   128 => x"84088105",
   129 => x"80dc840c",
   130 => x"80dc8408",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80dc84",
   134 => x"0c80dc80",
   135 => x"08810580",
   136 => x"dc800c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"dc880cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"dc880c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280dc",
   177 => x"88088407",
   178 => x"80dc880c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80d7",
   183 => x"f00c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80dc88",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80db",
   208 => x"f00c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02f8050d",
  1093 => x"80daac08",
  1094 => x"862a7083",
  1095 => x"068207e0",
  1096 => x"0c528051",
  1097 => x"86da2d86",
  1098 => x"c72d0288",
  1099 => x"050d0402",
  1100 => x"f8050d02",
  1101 => x"8f0580f5",
  1102 => x"2d80d7f8",
  1103 => x"08525270",
  1104 => x"80dd9d27",
  1105 => x"9a387171",
  1106 => x"81b72d80",
  1107 => x"d7f80881",
  1108 => x"0580d7f8",
  1109 => x"0c80d7f8",
  1110 => x"08518071",
  1111 => x"81b72d02",
  1112 => x"88050d04",
  1113 => x"02f4050d",
  1114 => x"7470842a",
  1115 => x"708f0680",
  1116 => x"d7f40805",
  1117 => x"7080f52d",
  1118 => x"54515353",
  1119 => x"a2af2d72",
  1120 => x"8f0680d7",
  1121 => x"f4080570",
  1122 => x"80f52d52",
  1123 => x"53a2af2d",
  1124 => x"028c050d",
  1125 => x"0402f405",
  1126 => x"0d747654",
  1127 => x"52727081",
  1128 => x"055480f5",
  1129 => x"2d517072",
  1130 => x"70810554",
  1131 => x"81b72d70",
  1132 => x"ec387072",
  1133 => x"81b72d02",
  1134 => x"8c050d04",
  1135 => x"02c4050d",
  1136 => x"800b80da",
  1137 => x"ac08a006",
  1138 => x"71725a40",
  1139 => x"405b810b",
  1140 => x"ec0c840b",
  1141 => x"ec0c6052",
  1142 => x"80dc8c51",
  1143 => x"80cb922d",
  1144 => x"80dbf008",
  1145 => x"7b2e8281",
  1146 => x"3880dc90",
  1147 => x"087bff12",
  1148 => x"575e5674",
  1149 => x"7b2e8b38",
  1150 => x"811d7581",
  1151 => x"2a565d74",
  1152 => x"f738f71d",
  1153 => x"5d815b80",
  1154 => x"762581dd",
  1155 => x"387c5274",
  1156 => x"5184a82d",
  1157 => x"80dde852",
  1158 => x"80dc8c51",
  1159 => x"80cde62d",
  1160 => x"80dbf008",
  1161 => x"802e81a7",
  1162 => x"3880dde8",
  1163 => x"5c83ff58",
  1164 => x"7e9c387b",
  1165 => x"7081055d",
  1166 => x"80f52d77",
  1167 => x"811959e4",
  1168 => x"0ce80cff",
  1169 => x"18587780",
  1170 => x"25e938a5",
  1171 => x"d7047b70",
  1172 => x"81055d80",
  1173 => x"f52d7781",
  1174 => x"1959e40c",
  1175 => x"f4800870",
  1176 => x"72327009",
  1177 => x"81057072",
  1178 => x"079f2a51",
  1179 => x"56565b59",
  1180 => x"7d80d038",
  1181 => x"81707406",
  1182 => x"54547280",
  1183 => x"2e80c438",
  1184 => x"7380dce0",
  1185 => x"0b80d7f8",
  1186 => x"0c80d688",
  1187 => x"5380dcdc",
  1188 => x"525ea395",
  1189 => x"2dff1770",
  1190 => x"5253a2e4",
  1191 => x"2d72882c",
  1192 => x"51a2e42d",
  1193 => x"a051a2af",
  1194 => x"2d7851a2",
  1195 => x"e42da051",
  1196 => x"a2af2d79",
  1197 => x"51a2e42d",
  1198 => x"80dcdc52",
  1199 => x"80dc9851",
  1200 => x"a3952dff",
  1201 => x"18587780",
  1202 => x"25ff8338",
  1203 => x"a5d70480",
  1204 => x"dbf0085b",
  1205 => x"84805680",
  1206 => x"dc8c5180",
  1207 => x"cdb52dfc",
  1208 => x"80168116",
  1209 => x"5656a487",
  1210 => x"0480dc90",
  1211 => x"08f80c7d",
  1212 => x"80d33880",
  1213 => x"d6537e84",
  1214 => x"3880cc53",
  1215 => x"7280dcdc",
  1216 => x"0b81b72d",
  1217 => x"80d69052",
  1218 => x"80dcdd51",
  1219 => x"a3952d80",
  1220 => x"dcdf0b80",
  1221 => x"d7f80c76",
  1222 => x"882c51a2",
  1223 => x"e42d7651",
  1224 => x"a2e42da0",
  1225 => x"51a2af2d",
  1226 => x"80dc9008",
  1227 => x"882a51a2",
  1228 => x"e42d80dc",
  1229 => x"900851a2",
  1230 => x"e42d80dc",
  1231 => x"dc5280dc",
  1232 => x"9851a395",
  1233 => x"2d805186",
  1234 => x"da2d7a80",
  1235 => x"2e883880",
  1236 => x"d7fc51a6",
  1237 => x"da0480d9",
  1238 => x"bc51afc1",
  1239 => x"2d7a80db",
  1240 => x"f00c02bc",
  1241 => x"050d0402",
  1242 => x"f0050d80",
  1243 => x"dcdc0b80",
  1244 => x"d7f80c80",
  1245 => x"0b80dcdc",
  1246 => x"0b81b72d",
  1247 => x"80d9e008",
  1248 => x"51a2e42d",
  1249 => x"ba51a2af",
  1250 => x"2d805480",
  1251 => x"d9e00814",
  1252 => x"e40cf480",
  1253 => x"0851a2e4",
  1254 => x"2da051a2",
  1255 => x"af2d8114",
  1256 => x"54877425",
  1257 => x"e63880dc",
  1258 => x"dc5280dc",
  1259 => x"9851a395",
  1260 => x"2d80d7fc",
  1261 => x"51afc12d",
  1262 => x"80d9e008",
  1263 => x"840580d9",
  1264 => x"e00c0290",
  1265 => x"050d0480",
  1266 => x"0b80d9e0",
  1267 => x"0c0402ec",
  1268 => x"050d840b",
  1269 => x"ec0cacfe",
  1270 => x"2da9b32d",
  1271 => x"81f92d83",
  1272 => x"53ace12d",
  1273 => x"8151858d",
  1274 => x"2dff1353",
  1275 => x"728025f1",
  1276 => x"38840bec",
  1277 => x"0c80d694",
  1278 => x"5186a02d",
  1279 => x"80c1bc2d",
  1280 => x"80dbf008",
  1281 => x"802e8194",
  1282 => x"38a3bc51",
  1283 => x"80d4bc2d",
  1284 => x"80d6ac52",
  1285 => x"80dc9851",
  1286 => x"a3952d80",
  1287 => x"d7fc51af",
  1288 => x"c12dada0",
  1289 => x"2da9bf2d",
  1290 => x"afd42d80",
  1291 => x"d8900b80",
  1292 => x"f52d80da",
  1293 => x"ac087081",
  1294 => x"06555654",
  1295 => x"72802e85",
  1296 => x"38738407",
  1297 => x"5474812a",
  1298 => x"70810651",
  1299 => x"5372802e",
  1300 => x"85387382",
  1301 => x"07547482",
  1302 => x"2a708106",
  1303 => x"51537280",
  1304 => x"2e853873",
  1305 => x"81075474",
  1306 => x"832a7081",
  1307 => x"06515372",
  1308 => x"802e8538",
  1309 => x"73880754",
  1310 => x"74842a70",
  1311 => x"81065153",
  1312 => x"72802e85",
  1313 => x"38739007",
  1314 => x"5473fc0c",
  1315 => x"865380db",
  1316 => x"f0088338",
  1317 => x"845372ec",
  1318 => x"0ca8a504",
  1319 => x"800b80db",
  1320 => x"f00c0294",
  1321 => x"050d0471",
  1322 => x"980c04ff",
  1323 => x"b00880db",
  1324 => x"f00c0481",
  1325 => x"0bffb00c",
  1326 => x"04800bff",
  1327 => x"b00c0402",
  1328 => x"f4050daa",
  1329 => x"cd0480db",
  1330 => x"f00881f0",
  1331 => x"2e098106",
  1332 => x"8a38810b",
  1333 => x"80daa40c",
  1334 => x"aacd0480",
  1335 => x"dbf00881",
  1336 => x"e02e0981",
  1337 => x"068a3881",
  1338 => x"0b80daa8",
  1339 => x"0caacd04",
  1340 => x"80dbf008",
  1341 => x"5280daa8",
  1342 => x"08802e89",
  1343 => x"3880dbf0",
  1344 => x"08818005",
  1345 => x"5271842c",
  1346 => x"728f0653",
  1347 => x"5380daa4",
  1348 => x"08802e9a",
  1349 => x"38728429",
  1350 => x"80d9e405",
  1351 => x"72138171",
  1352 => x"2b700973",
  1353 => x"0806730c",
  1354 => x"515353aa",
  1355 => x"c1047284",
  1356 => x"2980d9e4",
  1357 => x"05721383",
  1358 => x"712b7208",
  1359 => x"07720c53",
  1360 => x"53800b80",
  1361 => x"daa80c80",
  1362 => x"0b80daa4",
  1363 => x"0c80dda0",
  1364 => x"51abd42d",
  1365 => x"80dbf008",
  1366 => x"ff24feea",
  1367 => x"38800b80",
  1368 => x"dbf00c02",
  1369 => x"8c050d04",
  1370 => x"02f8050d",
  1371 => x"80d9e452",
  1372 => x"8f518072",
  1373 => x"70840554",
  1374 => x"0cff1151",
  1375 => x"708025f2",
  1376 => x"38028805",
  1377 => x"0d0402f0",
  1378 => x"050d7551",
  1379 => x"a9b92d70",
  1380 => x"822cfc06",
  1381 => x"80d9e411",
  1382 => x"72109e06",
  1383 => x"71087072",
  1384 => x"2a708306",
  1385 => x"82742b70",
  1386 => x"09740676",
  1387 => x"0c545156",
  1388 => x"57535153",
  1389 => x"a9b32d71",
  1390 => x"80dbf00c",
  1391 => x"0290050d",
  1392 => x"0402fc05",
  1393 => x"0d725180",
  1394 => x"710c800b",
  1395 => x"84120c02",
  1396 => x"84050d04",
  1397 => x"02f0050d",
  1398 => x"75700884",
  1399 => x"12085353",
  1400 => x"53ff5471",
  1401 => x"712ea838",
  1402 => x"a9b92d84",
  1403 => x"13087084",
  1404 => x"29148811",
  1405 => x"70087081",
  1406 => x"ff068418",
  1407 => x"08811187",
  1408 => x"06841a0c",
  1409 => x"53515551",
  1410 => x"5151a9b3",
  1411 => x"2d715473",
  1412 => x"80dbf00c",
  1413 => x"0290050d",
  1414 => x"0402f805",
  1415 => x"0da9b92d",
  1416 => x"e008708b",
  1417 => x"2a708106",
  1418 => x"51525270",
  1419 => x"802ea138",
  1420 => x"80dda008",
  1421 => x"70842980",
  1422 => x"dda80573",
  1423 => x"81ff0671",
  1424 => x"0c515180",
  1425 => x"dda00881",
  1426 => x"11870680",
  1427 => x"dda00c51",
  1428 => x"800b80dd",
  1429 => x"c80ca9ab",
  1430 => x"2da9b32d",
  1431 => x"0288050d",
  1432 => x"0402fc05",
  1433 => x"0da9b92d",
  1434 => x"810b80dd",
  1435 => x"c80ca9b3",
  1436 => x"2d80ddc8",
  1437 => x"085170f9",
  1438 => x"38028405",
  1439 => x"0d0402fc",
  1440 => x"050d80dd",
  1441 => x"a051abc1",
  1442 => x"2daae82d",
  1443 => x"ac9951a9",
  1444 => x"a72d0284",
  1445 => x"050d0480",
  1446 => x"ddd40880",
  1447 => x"dbf00c04",
  1448 => x"02fc050d",
  1449 => x"810b80da",
  1450 => x"b00c8151",
  1451 => x"858d2d02",
  1452 => x"84050d04",
  1453 => x"02fc050d",
  1454 => x"adbe04a9",
  1455 => x"bf2d80f6",
  1456 => x"51ab862d",
  1457 => x"80dbf008",
  1458 => x"f23880da",
  1459 => x"51ab862d",
  1460 => x"80dbf008",
  1461 => x"e63880db",
  1462 => x"f00880da",
  1463 => x"b00c80db",
  1464 => x"f0085185",
  1465 => x"8d2d0284",
  1466 => x"050d0402",
  1467 => x"ec050d76",
  1468 => x"54805287",
  1469 => x"0b881580",
  1470 => x"f52d5653",
  1471 => x"74722483",
  1472 => x"38a05372",
  1473 => x"5183842d",
  1474 => x"81128b15",
  1475 => x"80f52d54",
  1476 => x"52727225",
  1477 => x"de380294",
  1478 => x"050d0402",
  1479 => x"f0050d80",
  1480 => x"ddd40854",
  1481 => x"81f92d80",
  1482 => x"0b80ddd8",
  1483 => x"0c730880",
  1484 => x"2e818938",
  1485 => x"820b80dc",
  1486 => x"840c80dd",
  1487 => x"d8088f06",
  1488 => x"80dc800c",
  1489 => x"73085271",
  1490 => x"832e9638",
  1491 => x"71832689",
  1492 => x"3871812e",
  1493 => x"b038afa5",
  1494 => x"0471852e",
  1495 => x"a038afa5",
  1496 => x"04881480",
  1497 => x"f52d8415",
  1498 => x"0880d6bc",
  1499 => x"53545286",
  1500 => x"a02d7184",
  1501 => x"29137008",
  1502 => x"5252afa9",
  1503 => x"047351ad",
  1504 => x"eb2dafa5",
  1505 => x"0480daac",
  1506 => x"08881508",
  1507 => x"2c708106",
  1508 => x"51527180",
  1509 => x"2e883880",
  1510 => x"d6c051af",
  1511 => x"a20480d6",
  1512 => x"c45186a0",
  1513 => x"2d841408",
  1514 => x"5186a02d",
  1515 => x"80ddd808",
  1516 => x"810580dd",
  1517 => x"d80c8c14",
  1518 => x"54aead04",
  1519 => x"0290050d",
  1520 => x"047180dd",
  1521 => x"d40cae9b",
  1522 => x"2d80ddd8",
  1523 => x"08ff0580",
  1524 => x"dddc0c04",
  1525 => x"02e8050d",
  1526 => x"80ddd408",
  1527 => x"80dde008",
  1528 => x"575580f6",
  1529 => x"51ab862d",
  1530 => x"80dbf008",
  1531 => x"812a7081",
  1532 => x"06515271",
  1533 => x"802ea438",
  1534 => x"affe04a9",
  1535 => x"bf2d80f6",
  1536 => x"51ab862d",
  1537 => x"80dbf008",
  1538 => x"f23880da",
  1539 => x"b0088132",
  1540 => x"7080dab0",
  1541 => x"0c705252",
  1542 => x"858d2d80",
  1543 => x"0b80ddcc",
  1544 => x"0c800b80",
  1545 => x"ddd00c80",
  1546 => x"dab00883",
  1547 => x"8d3880da",
  1548 => x"51ab862d",
  1549 => x"80dbf008",
  1550 => x"802e8c38",
  1551 => x"80ddcc08",
  1552 => x"81800780",
  1553 => x"ddcc0c80",
  1554 => x"d951ab86",
  1555 => x"2d80dbf0",
  1556 => x"08802e8c",
  1557 => x"3880ddcc",
  1558 => x"0880c007",
  1559 => x"80ddcc0c",
  1560 => x"819451ab",
  1561 => x"862d80db",
  1562 => x"f008802e",
  1563 => x"8b3880dd",
  1564 => x"cc089007",
  1565 => x"80ddcc0c",
  1566 => x"819151ab",
  1567 => x"862d80db",
  1568 => x"f008802e",
  1569 => x"8b3880dd",
  1570 => x"cc08a007",
  1571 => x"80ddcc0c",
  1572 => x"81f551ab",
  1573 => x"862d80db",
  1574 => x"f008802e",
  1575 => x"8b3880dd",
  1576 => x"cc088107",
  1577 => x"80ddcc0c",
  1578 => x"81f251ab",
  1579 => x"862d80db",
  1580 => x"f008802e",
  1581 => x"8b3880dd",
  1582 => x"cc088207",
  1583 => x"80ddcc0c",
  1584 => x"81eb51ab",
  1585 => x"862d80db",
  1586 => x"f008802e",
  1587 => x"8b3880dd",
  1588 => x"cc088407",
  1589 => x"80ddcc0c",
  1590 => x"81f451ab",
  1591 => x"862d80db",
  1592 => x"f008802e",
  1593 => x"8b3880dd",
  1594 => x"cc088807",
  1595 => x"80ddcc0c",
  1596 => x"80d851ab",
  1597 => x"862d80db",
  1598 => x"f008802e",
  1599 => x"8c3880dd",
  1600 => x"d0088180",
  1601 => x"0780ddd0",
  1602 => x"0c9251ab",
  1603 => x"862d80db",
  1604 => x"f008802e",
  1605 => x"8c3880dd",
  1606 => x"d00880c0",
  1607 => x"0780ddd0",
  1608 => x"0c9451ab",
  1609 => x"862d80db",
  1610 => x"f008802e",
  1611 => x"8b3880dd",
  1612 => x"d0089007",
  1613 => x"80ddd00c",
  1614 => x"9151ab86",
  1615 => x"2d80dbf0",
  1616 => x"08802e8b",
  1617 => x"3880ddd0",
  1618 => x"08a00780",
  1619 => x"ddd00c9d",
  1620 => x"51ab862d",
  1621 => x"80dbf008",
  1622 => x"802e8b38",
  1623 => x"80ddd008",
  1624 => x"810780dd",
  1625 => x"d00c9b51",
  1626 => x"ab862d80",
  1627 => x"dbf00880",
  1628 => x"2e8b3880",
  1629 => x"ddd00882",
  1630 => x"0780ddd0",
  1631 => x"0c9c51ab",
  1632 => x"862d80db",
  1633 => x"f008802e",
  1634 => x"8b3880dd",
  1635 => x"d0088407",
  1636 => x"80ddd00c",
  1637 => x"a351ab86",
  1638 => x"2d80dbf0",
  1639 => x"08802e8b",
  1640 => x"3880ddd0",
  1641 => x"08880780",
  1642 => x"ddd00c81",
  1643 => x"fd51ab86",
  1644 => x"2d81fa51",
  1645 => x"ab862db9",
  1646 => x"8f0481f5",
  1647 => x"51ab862d",
  1648 => x"80dbf008",
  1649 => x"812a7081",
  1650 => x"06515271",
  1651 => x"802eb338",
  1652 => x"80dddc08",
  1653 => x"5271802e",
  1654 => x"8a38ff12",
  1655 => x"80dddc0c",
  1656 => x"b4820480",
  1657 => x"ddd80810",
  1658 => x"80ddd808",
  1659 => x"05708429",
  1660 => x"16515288",
  1661 => x"1208802e",
  1662 => x"8938ff51",
  1663 => x"88120852",
  1664 => x"712d81f2",
  1665 => x"51ab862d",
  1666 => x"80dbf008",
  1667 => x"812a7081",
  1668 => x"06515271",
  1669 => x"802eb438",
  1670 => x"80ddd808",
  1671 => x"ff1180dd",
  1672 => x"dc085653",
  1673 => x"53737225",
  1674 => x"8a388114",
  1675 => x"80dddc0c",
  1676 => x"b4cb0472",
  1677 => x"10137084",
  1678 => x"29165152",
  1679 => x"88120880",
  1680 => x"2e8938fe",
  1681 => x"51881208",
  1682 => x"52712d81",
  1683 => x"fd51ab86",
  1684 => x"2d80dbf0",
  1685 => x"08812a70",
  1686 => x"81065152",
  1687 => x"71802eb1",
  1688 => x"3880dddc",
  1689 => x"08802e8a",
  1690 => x"38800b80",
  1691 => x"dddc0cb5",
  1692 => x"910480dd",
  1693 => x"d8081080",
  1694 => x"ddd80805",
  1695 => x"70842916",
  1696 => x"51528812",
  1697 => x"08802e89",
  1698 => x"38fd5188",
  1699 => x"12085271",
  1700 => x"2d81fa51",
  1701 => x"ab862d80",
  1702 => x"dbf00881",
  1703 => x"2a708106",
  1704 => x"51527180",
  1705 => x"2eb13880",
  1706 => x"ddd808ff",
  1707 => x"11545280",
  1708 => x"dddc0873",
  1709 => x"25893872",
  1710 => x"80dddc0c",
  1711 => x"b5d70471",
  1712 => x"10127084",
  1713 => x"29165152",
  1714 => x"88120880",
  1715 => x"2e8938fc",
  1716 => x"51881208",
  1717 => x"52712d80",
  1718 => x"dddc0870",
  1719 => x"53547380",
  1720 => x"2e8a388c",
  1721 => x"15ff1555",
  1722 => x"55b5de04",
  1723 => x"820b80dc",
  1724 => x"840c718f",
  1725 => x"0680dc80",
  1726 => x"0c81eb51",
  1727 => x"ab862d80",
  1728 => x"dbf00881",
  1729 => x"2a708106",
  1730 => x"51527180",
  1731 => x"2ead3874",
  1732 => x"08852e09",
  1733 => x"8106a438",
  1734 => x"881580f5",
  1735 => x"2dff0552",
  1736 => x"71881681",
  1737 => x"b72d7198",
  1738 => x"2b527180",
  1739 => x"25883880",
  1740 => x"0b881681",
  1741 => x"b72d7451",
  1742 => x"adeb2d81",
  1743 => x"f451ab86",
  1744 => x"2d80dbf0",
  1745 => x"08812a70",
  1746 => x"81065152",
  1747 => x"71802eb3",
  1748 => x"38740885",
  1749 => x"2e098106",
  1750 => x"aa388815",
  1751 => x"80f52d81",
  1752 => x"05527188",
  1753 => x"1681b72d",
  1754 => x"7181ff06",
  1755 => x"8b1680f5",
  1756 => x"2d545272",
  1757 => x"72278738",
  1758 => x"72881681",
  1759 => x"b72d7451",
  1760 => x"adeb2d80",
  1761 => x"da51ab86",
  1762 => x"2d80dbf0",
  1763 => x"08812a70",
  1764 => x"81065152",
  1765 => x"71802e81",
  1766 => x"ad3880dd",
  1767 => x"d40880dd",
  1768 => x"dc085553",
  1769 => x"73802e8a",
  1770 => x"388c13ff",
  1771 => x"155553b7",
  1772 => x"a4047208",
  1773 => x"5271822e",
  1774 => x"a6387182",
  1775 => x"26893871",
  1776 => x"812eaa38",
  1777 => x"b8c60471",
  1778 => x"832eb438",
  1779 => x"71842e09",
  1780 => x"810680f2",
  1781 => x"38881308",
  1782 => x"51afc12d",
  1783 => x"b8c60480",
  1784 => x"dddc0851",
  1785 => x"88130852",
  1786 => x"712db8c6",
  1787 => x"04810b88",
  1788 => x"14082b80",
  1789 => x"daac0832",
  1790 => x"80daac0c",
  1791 => x"b89a0488",
  1792 => x"1380f52d",
  1793 => x"81058b14",
  1794 => x"80f52d53",
  1795 => x"54717424",
  1796 => x"83388054",
  1797 => x"73881481",
  1798 => x"b72dae9b",
  1799 => x"2db8c604",
  1800 => x"7508802e",
  1801 => x"a4387508",
  1802 => x"51ab862d",
  1803 => x"80dbf008",
  1804 => x"81065271",
  1805 => x"802e8c38",
  1806 => x"80dddc08",
  1807 => x"51841608",
  1808 => x"52712d88",
  1809 => x"165675d8",
  1810 => x"38805480",
  1811 => x"0b80dc84",
  1812 => x"0c738f06",
  1813 => x"80dc800c",
  1814 => x"a0527380",
  1815 => x"dddc082e",
  1816 => x"09810699",
  1817 => x"3880ddd8",
  1818 => x"08ff0574",
  1819 => x"32700981",
  1820 => x"05707207",
  1821 => x"9f2a9171",
  1822 => x"31515153",
  1823 => x"53715183",
  1824 => x"842d8114",
  1825 => x"548e7425",
  1826 => x"c23880da",
  1827 => x"b0085271",
  1828 => x"80dbf00c",
  1829 => x"0298050d",
  1830 => x"0402f405",
  1831 => x"0dd45281",
  1832 => x"ff720c71",
  1833 => x"085381ff",
  1834 => x"720c7288",
  1835 => x"2b83fe80",
  1836 => x"06720870",
  1837 => x"81ff0651",
  1838 => x"525381ff",
  1839 => x"720c7271",
  1840 => x"07882b72",
  1841 => x"087081ff",
  1842 => x"06515253",
  1843 => x"81ff720c",
  1844 => x"72710788",
  1845 => x"2b720870",
  1846 => x"81ff0672",
  1847 => x"0780dbf0",
  1848 => x"0c525302",
  1849 => x"8c050d04",
  1850 => x"02f4050d",
  1851 => x"74767181",
  1852 => x"ff06d40c",
  1853 => x"535380dd",
  1854 => x"e4088538",
  1855 => x"71892b52",
  1856 => x"71982ad4",
  1857 => x"0c71902a",
  1858 => x"7081ff06",
  1859 => x"d40c5171",
  1860 => x"882a7081",
  1861 => x"ff06d40c",
  1862 => x"517181ff",
  1863 => x"06d40c72",
  1864 => x"902a7081",
  1865 => x"ff06d40c",
  1866 => x"51d40870",
  1867 => x"81ff0651",
  1868 => x"5182b8bf",
  1869 => x"527081ff",
  1870 => x"2e098106",
  1871 => x"943881ff",
  1872 => x"0bd40cd4",
  1873 => x"087081ff",
  1874 => x"06ff1454",
  1875 => x"515171e5",
  1876 => x"387080db",
  1877 => x"f00c028c",
  1878 => x"050d0402",
  1879 => x"fc050d81",
  1880 => x"c75181ff",
  1881 => x"0bd40cff",
  1882 => x"11517080",
  1883 => x"25f43802",
  1884 => x"84050d04",
  1885 => x"02f4050d",
  1886 => x"81ff0bd4",
  1887 => x"0c935380",
  1888 => x"5287fc80",
  1889 => x"c151b9e8",
  1890 => x"2d80dbf0",
  1891 => x"088b3881",
  1892 => x"ff0bd40c",
  1893 => x"8153bba2",
  1894 => x"04badb2d",
  1895 => x"ff135372",
  1896 => x"de387280",
  1897 => x"dbf00c02",
  1898 => x"8c050d04",
  1899 => x"02ec050d",
  1900 => x"810b80dd",
  1901 => x"e40c8454",
  1902 => x"d008708f",
  1903 => x"2a708106",
  1904 => x"51515372",
  1905 => x"f33872d0",
  1906 => x"0cbadb2d",
  1907 => x"80d6c851",
  1908 => x"86a02dd0",
  1909 => x"08708f2a",
  1910 => x"70810651",
  1911 => x"515372f3",
  1912 => x"38810bd0",
  1913 => x"0cb15380",
  1914 => x"5284d480",
  1915 => x"c051b9e8",
  1916 => x"2d80dbf0",
  1917 => x"08812e93",
  1918 => x"3872822e",
  1919 => x"bf38ff13",
  1920 => x"5372e438",
  1921 => x"ff145473",
  1922 => x"ffae38ba",
  1923 => x"db2d83aa",
  1924 => x"52849c80",
  1925 => x"c851b9e8",
  1926 => x"2d80dbf0",
  1927 => x"08812e09",
  1928 => x"81069338",
  1929 => x"b9992d80",
  1930 => x"dbf00883",
  1931 => x"ffff0653",
  1932 => x"7283aa2e",
  1933 => x"9f38baf4",
  1934 => x"2dbccf04",
  1935 => x"80d6d451",
  1936 => x"86a02d80",
  1937 => x"53bea404",
  1938 => x"80d6ec51",
  1939 => x"86a02d80",
  1940 => x"54bdf504",
  1941 => x"81ff0bd4",
  1942 => x"0cb154ba",
  1943 => x"db2d8fcf",
  1944 => x"53805287",
  1945 => x"fc80f751",
  1946 => x"b9e82d80",
  1947 => x"dbf00855",
  1948 => x"80dbf008",
  1949 => x"812e0981",
  1950 => x"069c3881",
  1951 => x"ff0bd40c",
  1952 => x"820a5284",
  1953 => x"9c80e951",
  1954 => x"b9e82d80",
  1955 => x"dbf00880",
  1956 => x"2e8d38ba",
  1957 => x"db2dff13",
  1958 => x"5372c638",
  1959 => x"bde80481",
  1960 => x"ff0bd40c",
  1961 => x"80dbf008",
  1962 => x"5287fc80",
  1963 => x"fa51b9e8",
  1964 => x"2d80dbf0",
  1965 => x"08b23881",
  1966 => x"ff0bd40c",
  1967 => x"d4085381",
  1968 => x"ff0bd40c",
  1969 => x"81ff0bd4",
  1970 => x"0c81ff0b",
  1971 => x"d40c81ff",
  1972 => x"0bd40c72",
  1973 => x"862a7081",
  1974 => x"06765651",
  1975 => x"53729638",
  1976 => x"80dbf008",
  1977 => x"54bdf504",
  1978 => x"73822efe",
  1979 => x"db38ff14",
  1980 => x"5473fee7",
  1981 => x"387380dd",
  1982 => x"e40c738b",
  1983 => x"38815287",
  1984 => x"fc80d051",
  1985 => x"b9e82d81",
  1986 => x"ff0bd40c",
  1987 => x"d008708f",
  1988 => x"2a708106",
  1989 => x"51515372",
  1990 => x"f33872d0",
  1991 => x"0c81ff0b",
  1992 => x"d40c8153",
  1993 => x"7280dbf0",
  1994 => x"0c029405",
  1995 => x"0d0402e8",
  1996 => x"050d7855",
  1997 => x"805681ff",
  1998 => x"0bd40cd0",
  1999 => x"08708f2a",
  2000 => x"70810651",
  2001 => x"515372f3",
  2002 => x"3882810b",
  2003 => x"d00c81ff",
  2004 => x"0bd40c77",
  2005 => x"5287fc80",
  2006 => x"d151b9e8",
  2007 => x"2d80dbc6",
  2008 => x"df5480db",
  2009 => x"f008802e",
  2010 => x"8b3880d7",
  2011 => x"8c5186a0",
  2012 => x"2dbfc804",
  2013 => x"81ff0bd4",
  2014 => x"0cd40870",
  2015 => x"81ff0651",
  2016 => x"537281fe",
  2017 => x"2e098106",
  2018 => x"9e3880ff",
  2019 => x"53b9992d",
  2020 => x"80dbf008",
  2021 => x"75708405",
  2022 => x"570cff13",
  2023 => x"53728025",
  2024 => x"ec388156",
  2025 => x"bfad04ff",
  2026 => x"145473c8",
  2027 => x"3881ff0b",
  2028 => x"d40c81ff",
  2029 => x"0bd40cd0",
  2030 => x"08708f2a",
  2031 => x"70810651",
  2032 => x"515372f3",
  2033 => x"3872d00c",
  2034 => x"7580dbf0",
  2035 => x"0c029805",
  2036 => x"0d0402e8",
  2037 => x"050d7779",
  2038 => x"7b585555",
  2039 => x"80537276",
  2040 => x"25a43874",
  2041 => x"70810556",
  2042 => x"80f52d74",
  2043 => x"70810556",
  2044 => x"80f52d52",
  2045 => x"5271712e",
  2046 => x"87388151",
  2047 => x"80c08804",
  2048 => x"811353bf",
  2049 => x"de048051",
  2050 => x"7080dbf0",
  2051 => x"0c029805",
  2052 => x"0d0402ec",
  2053 => x"050d7655",
  2054 => x"74802e80",
  2055 => x"c4389a15",
  2056 => x"80e02d51",
  2057 => x"80cec02d",
  2058 => x"80dbf008",
  2059 => x"80dbf008",
  2060 => x"80e4980c",
  2061 => x"80dbf008",
  2062 => x"545480e3",
  2063 => x"f408802e",
  2064 => x"9b389415",
  2065 => x"80e02d51",
  2066 => x"80cec02d",
  2067 => x"80dbf008",
  2068 => x"902b83ff",
  2069 => x"f00a0670",
  2070 => x"75075153",
  2071 => x"7280e498",
  2072 => x"0c80e498",
  2073 => x"08537280",
  2074 => x"2e9e3880",
  2075 => x"e3ec08fe",
  2076 => x"14712980",
  2077 => x"e4800805",
  2078 => x"80e49c0c",
  2079 => x"70842b80",
  2080 => x"e3f80c54",
  2081 => x"80c1b704",
  2082 => x"80e48408",
  2083 => x"80e4980c",
  2084 => x"80e48808",
  2085 => x"80e49c0c",
  2086 => x"80e3f408",
  2087 => x"802e8c38",
  2088 => x"80e3ec08",
  2089 => x"842b5380",
  2090 => x"c1b20480",
  2091 => x"e48c0884",
  2092 => x"2b537280",
  2093 => x"e3f80c02",
  2094 => x"94050d04",
  2095 => x"02d8050d",
  2096 => x"800b80e3",
  2097 => x"f40c8454",
  2098 => x"bbac2d80",
  2099 => x"dbf00880",
  2100 => x"2e983880",
  2101 => x"dde85280",
  2102 => x"51beae2d",
  2103 => x"80dbf008",
  2104 => x"802e8738",
  2105 => x"fe5480c1",
  2106 => x"f204ff14",
  2107 => x"54738024",
  2108 => x"d738738e",
  2109 => x"3880d79c",
  2110 => x"5186a02d",
  2111 => x"735580c7",
  2112 => x"d0048056",
  2113 => x"810b80e4",
  2114 => x"a00c8853",
  2115 => x"80d7b052",
  2116 => x"80de9e51",
  2117 => x"bfd22d80",
  2118 => x"dbf00876",
  2119 => x"2e098106",
  2120 => x"893880db",
  2121 => x"f00880e4",
  2122 => x"a00c8853",
  2123 => x"80d7bc52",
  2124 => x"80deba51",
  2125 => x"bfd22d80",
  2126 => x"dbf00889",
  2127 => x"3880dbf0",
  2128 => x"0880e4a0",
  2129 => x"0c80e4a0",
  2130 => x"08802e81",
  2131 => x"843880e1",
  2132 => x"ae0b80f5",
  2133 => x"2d80e1af",
  2134 => x"0b80f52d",
  2135 => x"71982b71",
  2136 => x"902b0780",
  2137 => x"e1b00b80",
  2138 => x"f52d7088",
  2139 => x"2b720780",
  2140 => x"e1b10b80",
  2141 => x"f52d7107",
  2142 => x"80e1e60b",
  2143 => x"80f52d80",
  2144 => x"e1e70b80",
  2145 => x"f52d7188",
  2146 => x"2b07535f",
  2147 => x"54525a56",
  2148 => x"57557381",
  2149 => x"abaa2e09",
  2150 => x"81069038",
  2151 => x"755180ce",
  2152 => x"8f2d80db",
  2153 => x"f0085680",
  2154 => x"c3ba0473",
  2155 => x"82d4d52e",
  2156 => x"893880d7",
  2157 => x"c85180c4",
  2158 => x"870480dd",
  2159 => x"e8527551",
  2160 => x"beae2d80",
  2161 => x"dbf00855",
  2162 => x"80dbf008",
  2163 => x"802e8480",
  2164 => x"38885380",
  2165 => x"d7bc5280",
  2166 => x"deba51bf",
  2167 => x"d22d80db",
  2168 => x"f0088b38",
  2169 => x"810b80e3",
  2170 => x"f40c80c4",
  2171 => x"8e048853",
  2172 => x"80d7b052",
  2173 => x"80de9e51",
  2174 => x"bfd22d80",
  2175 => x"dbf00880",
  2176 => x"2e8c3880",
  2177 => x"d7dc5186",
  2178 => x"a02d80c4",
  2179 => x"ed0480e1",
  2180 => x"e60b80f5",
  2181 => x"2d547380",
  2182 => x"d52e0981",
  2183 => x"0680ce38",
  2184 => x"80e1e70b",
  2185 => x"80f52d54",
  2186 => x"7381aa2e",
  2187 => x"098106bd",
  2188 => x"38800b80",
  2189 => x"dde80b80",
  2190 => x"f52d5654",
  2191 => x"7481e92e",
  2192 => x"83388154",
  2193 => x"7481eb2e",
  2194 => x"8c388055",
  2195 => x"73752e09",
  2196 => x"810682fc",
  2197 => x"3880ddf3",
  2198 => x"0b80f52d",
  2199 => x"55748e38",
  2200 => x"80ddf40b",
  2201 => x"80f52d54",
  2202 => x"73822e87",
  2203 => x"38805580",
  2204 => x"c7d00480",
  2205 => x"ddf50b80",
  2206 => x"f52d7080",
  2207 => x"e3ec0cff",
  2208 => x"0580e3f0",
  2209 => x"0c80ddf6",
  2210 => x"0b80f52d",
  2211 => x"80ddf70b",
  2212 => x"80f52d58",
  2213 => x"76057782",
  2214 => x"80290570",
  2215 => x"80e3fc0c",
  2216 => x"80ddf80b",
  2217 => x"80f52d70",
  2218 => x"80e4900c",
  2219 => x"80e3f408",
  2220 => x"59575876",
  2221 => x"802e81b8",
  2222 => x"38885380",
  2223 => x"d7bc5280",
  2224 => x"deba51bf",
  2225 => x"d22d80db",
  2226 => x"f0088284",
  2227 => x"3880e3ec",
  2228 => x"0870842b",
  2229 => x"80e3f80c",
  2230 => x"7080e48c",
  2231 => x"0c80de8d",
  2232 => x"0b80f52d",
  2233 => x"80de8c0b",
  2234 => x"80f52d71",
  2235 => x"82802905",
  2236 => x"80de8e0b",
  2237 => x"80f52d70",
  2238 => x"84808029",
  2239 => x"1280de8f",
  2240 => x"0b80f52d",
  2241 => x"7081800a",
  2242 => x"29127080",
  2243 => x"e4940c80",
  2244 => x"e4900871",
  2245 => x"2980e3fc",
  2246 => x"08057080",
  2247 => x"e4800c80",
  2248 => x"de950b80",
  2249 => x"f52d80de",
  2250 => x"940b80f5",
  2251 => x"2d718280",
  2252 => x"290580de",
  2253 => x"960b80f5",
  2254 => x"2d708480",
  2255 => x"80291280",
  2256 => x"de970b80",
  2257 => x"f52d7098",
  2258 => x"2b81f00a",
  2259 => x"06720570",
  2260 => x"80e4840c",
  2261 => x"fe117e29",
  2262 => x"770580e4",
  2263 => x"880c5259",
  2264 => x"5243545e",
  2265 => x"51525952",
  2266 => x"5d575957",
  2267 => x"80c7c804",
  2268 => x"80ddfa0b",
  2269 => x"80f52d80",
  2270 => x"ddf90b80",
  2271 => x"f52d7182",
  2272 => x"80290570",
  2273 => x"80e3f80c",
  2274 => x"70a02983",
  2275 => x"ff057089",
  2276 => x"2a7080e4",
  2277 => x"8c0c80dd",
  2278 => x"ff0b80f5",
  2279 => x"2d80ddfe",
  2280 => x"0b80f52d",
  2281 => x"71828029",
  2282 => x"057080e4",
  2283 => x"940c7b71",
  2284 => x"291e7080",
  2285 => x"e4880c7d",
  2286 => x"80e4840c",
  2287 => x"730580e4",
  2288 => x"800c555e",
  2289 => x"51515555",
  2290 => x"805180c0",
  2291 => x"922d8155",
  2292 => x"7480dbf0",
  2293 => x"0c02a805",
  2294 => x"0d0402ec",
  2295 => x"050d7670",
  2296 => x"872c7180",
  2297 => x"ff065556",
  2298 => x"5480e3f4",
  2299 => x"088a3873",
  2300 => x"882c7481",
  2301 => x"ff065455",
  2302 => x"80dde852",
  2303 => x"80e3fc08",
  2304 => x"1551beae",
  2305 => x"2d80dbf0",
  2306 => x"085480db",
  2307 => x"f008802e",
  2308 => x"bb3880e3",
  2309 => x"f408802e",
  2310 => x"9c387284",
  2311 => x"2980dde8",
  2312 => x"05700852",
  2313 => x"5380ce8f",
  2314 => x"2d80dbf0",
  2315 => x"08f00a06",
  2316 => x"5380c8ca",
  2317 => x"04721080",
  2318 => x"dde80570",
  2319 => x"80e02d52",
  2320 => x"5380cec0",
  2321 => x"2d80dbf0",
  2322 => x"08537254",
  2323 => x"7380dbf0",
  2324 => x"0c029405",
  2325 => x"0d0402e0",
  2326 => x"050d7970",
  2327 => x"842c80e4",
  2328 => x"9c080571",
  2329 => x"8f065255",
  2330 => x"53728a38",
  2331 => x"80dde852",
  2332 => x"7351beae",
  2333 => x"2d72a029",
  2334 => x"80dde805",
  2335 => x"54807480",
  2336 => x"f52d5653",
  2337 => x"74732e83",
  2338 => x"38815374",
  2339 => x"81e52e81",
  2340 => x"f5388170",
  2341 => x"74065458",
  2342 => x"72802e81",
  2343 => x"e9388b14",
  2344 => x"80f52d70",
  2345 => x"832a7906",
  2346 => x"5856769c",
  2347 => x"3880dab4",
  2348 => x"08537289",
  2349 => x"387280e1",
  2350 => x"e80b81b7",
  2351 => x"2d7680da",
  2352 => x"b40c7353",
  2353 => x"80cb8804",
  2354 => x"758f2e09",
  2355 => x"810681b6",
  2356 => x"38749f06",
  2357 => x"8d2980e1",
  2358 => x"db115153",
  2359 => x"811480f5",
  2360 => x"2d737081",
  2361 => x"055581b7",
  2362 => x"2d831480",
  2363 => x"f52d7370",
  2364 => x"81055581",
  2365 => x"b72d8514",
  2366 => x"80f52d73",
  2367 => x"70810555",
  2368 => x"81b72d87",
  2369 => x"1480f52d",
  2370 => x"73708105",
  2371 => x"5581b72d",
  2372 => x"891480f5",
  2373 => x"2d737081",
  2374 => x"055581b7",
  2375 => x"2d8e1480",
  2376 => x"f52d7370",
  2377 => x"81055581",
  2378 => x"b72d9014",
  2379 => x"80f52d73",
  2380 => x"70810555",
  2381 => x"81b72d92",
  2382 => x"1480f52d",
  2383 => x"73708105",
  2384 => x"5581b72d",
  2385 => x"941480f5",
  2386 => x"2d737081",
  2387 => x"055581b7",
  2388 => x"2d961480",
  2389 => x"f52d7370",
  2390 => x"81055581",
  2391 => x"b72d9814",
  2392 => x"80f52d73",
  2393 => x"70810555",
  2394 => x"81b72d9c",
  2395 => x"1480f52d",
  2396 => x"73708105",
  2397 => x"5581b72d",
  2398 => x"9e1480f5",
  2399 => x"2d7381b7",
  2400 => x"2d7780da",
  2401 => x"b40c8053",
  2402 => x"7280dbf0",
  2403 => x"0c02a005",
  2404 => x"0d0402cc",
  2405 => x"050d7e60",
  2406 => x"5e5a800b",
  2407 => x"80e49808",
  2408 => x"80e49c08",
  2409 => x"595c5680",
  2410 => x"5880e3f8",
  2411 => x"08782e81",
  2412 => x"bc38778f",
  2413 => x"06a01757",
  2414 => x"54739138",
  2415 => x"80dde852",
  2416 => x"76518117",
  2417 => x"57beae2d",
  2418 => x"80dde856",
  2419 => x"807680f5",
  2420 => x"2d565474",
  2421 => x"742e8338",
  2422 => x"81547481",
  2423 => x"e52e8181",
  2424 => x"38817075",
  2425 => x"06555c73",
  2426 => x"802e80f5",
  2427 => x"388b1680",
  2428 => x"f52d9806",
  2429 => x"597880e9",
  2430 => x"388b537c",
  2431 => x"527551bf",
  2432 => x"d22d80db",
  2433 => x"f00880d9",
  2434 => x"389c1608",
  2435 => x"5180ce8f",
  2436 => x"2d80dbf0",
  2437 => x"08841b0c",
  2438 => x"9a1680e0",
  2439 => x"2d5180ce",
  2440 => x"c02d80db",
  2441 => x"f00880db",
  2442 => x"f008881c",
  2443 => x"0c80dbf0",
  2444 => x"08555580",
  2445 => x"e3f40880",
  2446 => x"2e9a3894",
  2447 => x"1680e02d",
  2448 => x"5180cec0",
  2449 => x"2d80dbf0",
  2450 => x"08902b83",
  2451 => x"fff00a06",
  2452 => x"70165154",
  2453 => x"73881b0c",
  2454 => x"787a0c7b",
  2455 => x"5480cdab",
  2456 => x"04811858",
  2457 => x"80e3f808",
  2458 => x"7826fec6",
  2459 => x"3880e3f4",
  2460 => x"08802eb5",
  2461 => x"387a5180",
  2462 => x"c7da2d80",
  2463 => x"dbf00880",
  2464 => x"dbf00880",
  2465 => x"fffffff8",
  2466 => x"06555b73",
  2467 => x"80ffffff",
  2468 => x"f82e9638",
  2469 => x"80dbf008",
  2470 => x"fe0580e3",
  2471 => x"ec082980",
  2472 => x"e4800805",
  2473 => x"5780cba7",
  2474 => x"04805473",
  2475 => x"80dbf00c",
  2476 => x"02b4050d",
  2477 => x"0402f405",
  2478 => x"0d747008",
  2479 => x"8105710c",
  2480 => x"700880e3",
  2481 => x"f0080653",
  2482 => x"53719038",
  2483 => x"88130851",
  2484 => x"80c7da2d",
  2485 => x"80dbf008",
  2486 => x"88140c81",
  2487 => x"0b80dbf0",
  2488 => x"0c028c05",
  2489 => x"0d0402f0",
  2490 => x"050d7588",
  2491 => x"1108fe05",
  2492 => x"80e3ec08",
  2493 => x"2980e480",
  2494 => x"08117208",
  2495 => x"80e3f008",
  2496 => x"06057955",
  2497 => x"535454be",
  2498 => x"ae2d0290",
  2499 => x"050d0402",
  2500 => x"f4050d74",
  2501 => x"70882a83",
  2502 => x"fe800670",
  2503 => x"72982a07",
  2504 => x"72882b87",
  2505 => x"fc808006",
  2506 => x"73982b81",
  2507 => x"f00a0671",
  2508 => x"73070780",
  2509 => x"dbf00c56",
  2510 => x"51535102",
  2511 => x"8c050d04",
  2512 => x"02f8050d",
  2513 => x"028e0580",
  2514 => x"f52d7488",
  2515 => x"2b077083",
  2516 => x"ffff0680",
  2517 => x"dbf00c51",
  2518 => x"0288050d",
  2519 => x"0402f405",
  2520 => x"0d747678",
  2521 => x"53545280",
  2522 => x"71259738",
  2523 => x"72708105",
  2524 => x"5480f52d",
  2525 => x"72708105",
  2526 => x"5481b72d",
  2527 => x"ff115170",
  2528 => x"eb388072",
  2529 => x"81b72d02",
  2530 => x"8c050d04",
  2531 => x"02e8050d",
  2532 => x"77568070",
  2533 => x"56547376",
  2534 => x"24b73880",
  2535 => x"e3f80874",
  2536 => x"2eaf3873",
  2537 => x"5180c8d6",
  2538 => x"2d80dbf0",
  2539 => x"0880dbf0",
  2540 => x"08098105",
  2541 => x"7080dbf0",
  2542 => x"08079f2a",
  2543 => x"77058117",
  2544 => x"57575353",
  2545 => x"74762489",
  2546 => x"3880e3f8",
  2547 => x"087426d3",
  2548 => x"387280db",
  2549 => x"f00c0298",
  2550 => x"050d0402",
  2551 => x"f0050d80",
  2552 => x"dbec0816",
  2553 => x"5180cf8c",
  2554 => x"2d80dbf0",
  2555 => x"08802ea0",
  2556 => x"388b5380",
  2557 => x"dbf00852",
  2558 => x"80e1e851",
  2559 => x"80cedd2d",
  2560 => x"80e4a408",
  2561 => x"5473802e",
  2562 => x"873880e1",
  2563 => x"e851732d",
  2564 => x"0290050d",
  2565 => x"0402dc05",
  2566 => x"0d80705a",
  2567 => x"557480db",
  2568 => x"ec0825b5",
  2569 => x"3880e3f8",
  2570 => x"08752ead",
  2571 => x"38785180",
  2572 => x"c8d62d80",
  2573 => x"dbf00809",
  2574 => x"81057080",
  2575 => x"dbf00807",
  2576 => x"9f2a7605",
  2577 => x"811b5b56",
  2578 => x"547480db",
  2579 => x"ec082589",
  2580 => x"3880e3f8",
  2581 => x"087926d5",
  2582 => x"38805578",
  2583 => x"80e3f808",
  2584 => x"2781e438",
  2585 => x"785180c8",
  2586 => x"d62d80db",
  2587 => x"f008802e",
  2588 => x"81b43880",
  2589 => x"dbf0088b",
  2590 => x"0580f52d",
  2591 => x"70842a70",
  2592 => x"81067710",
  2593 => x"78842b80",
  2594 => x"e1e80b80",
  2595 => x"f52d5c5c",
  2596 => x"53515556",
  2597 => x"73802e80",
  2598 => x"ce387416",
  2599 => x"822b80d2",
  2600 => x"eb0b80da",
  2601 => x"c0120c54",
  2602 => x"77753110",
  2603 => x"80e4a811",
  2604 => x"55569074",
  2605 => x"70810556",
  2606 => x"81b72da0",
  2607 => x"7481b72d",
  2608 => x"7681ff06",
  2609 => x"81165854",
  2610 => x"73802e8b",
  2611 => x"389c5380",
  2612 => x"e1e85280",
  2613 => x"d1de048b",
  2614 => x"5380dbf0",
  2615 => x"085280e4",
  2616 => x"aa165180",
  2617 => x"d29c0474",
  2618 => x"16822b80",
  2619 => x"cfdb0b80",
  2620 => x"dac0120c",
  2621 => x"547681ff",
  2622 => x"06811658",
  2623 => x"5473802e",
  2624 => x"8b389c53",
  2625 => x"80e1e852",
  2626 => x"80d29304",
  2627 => x"8b5380db",
  2628 => x"f0085277",
  2629 => x"75311080",
  2630 => x"e4a80551",
  2631 => x"765580ce",
  2632 => x"dd2d80d2",
  2633 => x"bb047490",
  2634 => x"29753170",
  2635 => x"1080e4a8",
  2636 => x"05515480",
  2637 => x"dbf00874",
  2638 => x"81b72d81",
  2639 => x"1959748b",
  2640 => x"24a43880",
  2641 => x"d0db0474",
  2642 => x"90297531",
  2643 => x"701080e4",
  2644 => x"a8058c77",
  2645 => x"31575154",
  2646 => x"807481b7",
  2647 => x"2d9e14ff",
  2648 => x"16565474",
  2649 => x"f33802a4",
  2650 => x"050d0402",
  2651 => x"fc050d80",
  2652 => x"dbec0813",
  2653 => x"5180cf8c",
  2654 => x"2d80dbf0",
  2655 => x"08802e8a",
  2656 => x"3880dbf0",
  2657 => x"085180c0",
  2658 => x"922d800b",
  2659 => x"80dbec0c",
  2660 => x"80d0952d",
  2661 => x"ae9b2d02",
  2662 => x"84050d04",
  2663 => x"02fc050d",
  2664 => x"725170fd",
  2665 => x"2eb23870",
  2666 => x"fd248b38",
  2667 => x"70fc2e80",
  2668 => x"d03880d4",
  2669 => x"8b0470fe",
  2670 => x"2eb93870",
  2671 => x"ff2e0981",
  2672 => x"0680c838",
  2673 => x"80dbec08",
  2674 => x"5170802e",
  2675 => x"be38ff11",
  2676 => x"80dbec0c",
  2677 => x"80d48b04",
  2678 => x"80dbec08",
  2679 => x"f0057080",
  2680 => x"dbec0c51",
  2681 => x"708025a3",
  2682 => x"38800b80",
  2683 => x"dbec0c80",
  2684 => x"d48b0480",
  2685 => x"dbec0881",
  2686 => x"0580dbec",
  2687 => x"0c80d48b",
  2688 => x"0480dbec",
  2689 => x"08900580",
  2690 => x"dbec0c80",
  2691 => x"d0952dae",
  2692 => x"9b2d0284",
  2693 => x"050d0402",
  2694 => x"fc050d80",
  2695 => x"0b80dbec",
  2696 => x"0c80d095",
  2697 => x"2dad972d",
  2698 => x"80dbf008",
  2699 => x"80dbdc0c",
  2700 => x"80dab851",
  2701 => x"afc12d02",
  2702 => x"84050d04",
  2703 => x"7180e4a4",
  2704 => x"0c040000",
  2705 => x"00ffffff",
  2706 => x"ff00ffff",
  2707 => x"ffff00ff",
  2708 => x"ffffff00",
  2709 => x"30313233",
  2710 => x"34353637",
  2711 => x"38394142",
  2712 => x"43444546",
  2713 => x"00000000",
  2714 => x"44656275",
  2715 => x"67000000",
  2716 => x"52657365",
  2717 => x"74000000",
  2718 => x"5363616e",
  2719 => x"6c696e65",
  2720 => x"73000000",
  2721 => x"50414c20",
  2722 => x"2f204e54",
  2723 => x"53430000",
  2724 => x"436f6c6f",
  2725 => x"72000000",
  2726 => x"44696666",
  2727 => x"6963756c",
  2728 => x"74792041",
  2729 => x"00000000",
  2730 => x"44696666",
  2731 => x"6963756c",
  2732 => x"74792042",
  2733 => x"00000000",
  2734 => x"56657269",
  2735 => x"66790000",
  2736 => x"524f4d00",
  2737 => x"626f6f74",
  2738 => x"00000000",
  2739 => x"53656c65",
  2740 => x"63740000",
  2741 => x"53746172",
  2742 => x"74000000",
  2743 => x"4c6f6164",
  2744 => x"20524f4d",
  2745 => x"20100000",
  2746 => x"45786974",
  2747 => x"00000000",
  2748 => x"524f4d20",
  2749 => x"6c6f6164",
  2750 => x"696e6720",
  2751 => x"6661696c",
  2752 => x"65640000",
  2753 => x"4f4b0000",
  2754 => x"45525220",
  2755 => x"00000000",
  2756 => x"4f4b2000",
  2757 => x"496e6974",
  2758 => x"69616c69",
  2759 => x"7a696e67",
  2760 => x"20534420",
  2761 => x"63617264",
  2762 => x"0a000000",
  2763 => x"436f6c6c",
  2764 => x"6563746f",
  2765 => x"72566973",
  2766 => x"696f6e00",
  2767 => x"16200000",
  2768 => x"14200000",
  2769 => x"15200000",
  2770 => x"53442069",
  2771 => x"6e69742e",
  2772 => x"2e2e0a00",
  2773 => x"53442063",
  2774 => x"61726420",
  2775 => x"72657365",
  2776 => x"74206661",
  2777 => x"696c6564",
  2778 => x"210a0000",
  2779 => x"53444843",
  2780 => x"20657272",
  2781 => x"6f72210a",
  2782 => x"00000000",
  2783 => x"57726974",
  2784 => x"65206661",
  2785 => x"696c6564",
  2786 => x"0a000000",
  2787 => x"52656164",
  2788 => x"20666169",
  2789 => x"6c65640a",
  2790 => x"00000000",
  2791 => x"43617264",
  2792 => x"20696e69",
  2793 => x"74206661",
  2794 => x"696c6564",
  2795 => x"0a000000",
  2796 => x"46415431",
  2797 => x"36202020",
  2798 => x"00000000",
  2799 => x"46415433",
  2800 => x"32202020",
  2801 => x"00000000",
  2802 => x"4e6f2070",
  2803 => x"61727469",
  2804 => x"74696f6e",
  2805 => x"20736967",
  2806 => x"0a000000",
  2807 => x"42616420",
  2808 => x"70617274",
  2809 => x"0a000000",
  2810 => x"4261636b",
  2811 => x"00000000",
  2812 => x"00000002",
  2813 => x"00002a54",
  2814 => x"00002e5c",
  2815 => x"00000002",
  2816 => x"00002e18",
  2817 => x"000013c7",
  2818 => x"00000002",
  2819 => x"00002a68",
  2820 => x"00001367",
  2821 => x"00000002",
  2822 => x"00002a70",
  2823 => x"0000035a",
  2824 => x"00000001",
  2825 => x"00002a78",
  2826 => x"00000000",
  2827 => x"00000001",
  2828 => x"00002a84",
  2829 => x"00000001",
  2830 => x"00000001",
  2831 => x"00002a90",
  2832 => x"00000002",
  2833 => x"00000001",
  2834 => x"00002a98",
  2835 => x"00000003",
  2836 => x"00000001",
  2837 => x"00002aa8",
  2838 => x"00000004",
  2839 => x"00000001",
  2840 => x"00002ab8",
  2841 => x"00000005",
  2842 => x"00000001",
  2843 => x"00002ac0",
  2844 => x"00000006",
  2845 => x"00000002",
  2846 => x"00002ac4",
  2847 => x"00001110",
  2848 => x"00000002",
  2849 => x"00002acc",
  2850 => x"0000036e",
  2851 => x"00000002",
  2852 => x"00002ad4",
  2853 => x"00000a3f",
  2854 => x"00000002",
  2855 => x"00002adc",
  2856 => x"00002a17",
  2857 => x"00000002",
  2858 => x"00002ae8",
  2859 => x"000016b4",
  2860 => x"00000000",
  2861 => x"00000000",
  2862 => x"00000000",
  2863 => x"00000004",
  2864 => x"00002af0",
  2865 => x"00002cbc",
  2866 => x"00000004",
  2867 => x"00002b04",
  2868 => x"00002bfc",
  2869 => x"00000000",
  2870 => x"00000000",
  2871 => x"00000000",
  2872 => x"00000000",
  2873 => x"00000000",
  2874 => x"00000000",
  2875 => x"00000000",
  2876 => x"00000000",
  2877 => x"00000000",
  2878 => x"00000000",
  2879 => x"00000000",
  2880 => x"00000000",
  2881 => x"00000000",
  2882 => x"00000000",
  2883 => x"00000000",
  2884 => x"00000000",
  2885 => x"00000000",
  2886 => x"00000000",
  2887 => x"00000000",
  2888 => x"00000000",
  2889 => x"00000000",
  2890 => x"00000000",
  2891 => x"00000006",
  2892 => x"00000000",
  2893 => x"00000000",
  2894 => x"00000002",
  2895 => x"00003228",
  2896 => x"000027db",
  2897 => x"00000002",
  2898 => x"00003246",
  2899 => x"000027db",
  2900 => x"00000002",
  2901 => x"00003264",
  2902 => x"000027db",
  2903 => x"00000002",
  2904 => x"00003282",
  2905 => x"000027db",
  2906 => x"00000002",
  2907 => x"000032a0",
  2908 => x"000027db",
  2909 => x"00000002",
  2910 => x"000032be",
  2911 => x"000027db",
  2912 => x"00000002",
  2913 => x"000032dc",
  2914 => x"000027db",
  2915 => x"00000002",
  2916 => x"000032fa",
  2917 => x"000027db",
  2918 => x"00000002",
  2919 => x"00003318",
  2920 => x"000027db",
  2921 => x"00000002",
  2922 => x"00003336",
  2923 => x"000027db",
  2924 => x"00000002",
  2925 => x"00003354",
  2926 => x"000027db",
  2927 => x"00000002",
  2928 => x"00003372",
  2929 => x"000027db",
  2930 => x"00000002",
  2931 => x"00003390",
  2932 => x"000027db",
  2933 => x"00000004",
  2934 => x"00002be8",
  2935 => x"00000000",
  2936 => x"00000000",
  2937 => x"00000000",
  2938 => x"0000299c",
  2939 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

