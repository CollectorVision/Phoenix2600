-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80db",
     9 => x"e0080b0b",
    10 => x"80dbe408",
    11 => x"0b0b80db",
    12 => x"e8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"dbe80c0b",
    16 => x"0b80dbe4",
    17 => x"0c0b0b80",
    18 => x"dbe00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d4bc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80dbe070",
    57 => x"80e7a027",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a5e6",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80db",
    65 => x"f00c9f0b",
    66 => x"80dbf40c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"dbf408ff",
    70 => x"0580dbf4",
    71 => x"0c80dbf4",
    72 => x"088025e8",
    73 => x"3880dbf0",
    74 => x"08ff0580",
    75 => x"dbf00c80",
    76 => x"dbf00880",
    77 => x"25d03880",
    78 => x"0b80dbf4",
    79 => x"0c800b80",
    80 => x"dbf00c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80dbf008",
   100 => x"25913882",
   101 => x"c82d80db",
   102 => x"f008ff05",
   103 => x"80dbf00c",
   104 => x"838a0480",
   105 => x"dbf00880",
   106 => x"dbf40853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80dbf008",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"dbf40881",
   116 => x"0580dbf4",
   117 => x"0c80dbf4",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80dbf4",
   121 => x"0c80dbf0",
   122 => x"08810580",
   123 => x"dbf00c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480db",
   128 => x"f4088105",
   129 => x"80dbf40c",
   130 => x"80dbf408",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80dbf4",
   134 => x"0c80dbf0",
   135 => x"08810580",
   136 => x"dbf00c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"dbf80cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"dbf80c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280db",
   177 => x"f8088407",
   178 => x"80dbf80c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80d7",
   183 => x"e00c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80dbf8",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80db",
   208 => x"e00c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02f8050d",
  1093 => x"028f0580",
  1094 => x"f52d80d7",
  1095 => x"e8085252",
  1096 => x"7080dd8d",
  1097 => x"279a3871",
  1098 => x"7181b72d",
  1099 => x"80d7e808",
  1100 => x"810580d7",
  1101 => x"e80c80d7",
  1102 => x"e8085180",
  1103 => x"7181b72d",
  1104 => x"0288050d",
  1105 => x"0402f405",
  1106 => x"0d747084",
  1107 => x"2a708f06",
  1108 => x"80d7e408",
  1109 => x"057080f5",
  1110 => x"2d545153",
  1111 => x"53a2902d",
  1112 => x"728f0680",
  1113 => x"d7e40805",
  1114 => x"7080f52d",
  1115 => x"5253a290",
  1116 => x"2d028c05",
  1117 => x"0d0402f4",
  1118 => x"050d7476",
  1119 => x"54527270",
  1120 => x"81055480",
  1121 => x"f52d5170",
  1122 => x"72708105",
  1123 => x"5481b72d",
  1124 => x"70ec3870",
  1125 => x"7281b72d",
  1126 => x"028c050d",
  1127 => x"0402d005",
  1128 => x"0d800b80",
  1129 => x"da9c0881",
  1130 => x"8006715d",
  1131 => x"5d59810b",
  1132 => x"ec0c840b",
  1133 => x"ec0c7d52",
  1134 => x"80dbfc51",
  1135 => x"80cb8a2d",
  1136 => x"80dbe008",
  1137 => x"792e80ff",
  1138 => x"3880dc80",
  1139 => x"0879ff12",
  1140 => x"57595774",
  1141 => x"792e8b38",
  1142 => x"81187581",
  1143 => x"2a565874",
  1144 => x"f738f718",
  1145 => x"58815980",
  1146 => x"772580db",
  1147 => x"38775274",
  1148 => x"5184a82d",
  1149 => x"80ddd852",
  1150 => x"80dbfc51",
  1151 => x"80cdde2d",
  1152 => x"80dbe008",
  1153 => x"802ea638",
  1154 => x"80ddd85a",
  1155 => x"7ba73883",
  1156 => x"ff567970",
  1157 => x"81055b80",
  1158 => x"f52d7b81",
  1159 => x"1d5de40c",
  1160 => x"e80cff16",
  1161 => x"56758025",
  1162 => x"e938a4b5",
  1163 => x"0480dbe0",
  1164 => x"08598480",
  1165 => x"5780dbfc",
  1166 => x"5180cdad",
  1167 => x"2dfc8017",
  1168 => x"81165657",
  1169 => x"a3e70480",
  1170 => x"dc8008f8",
  1171 => x"0c810be0",
  1172 => x"0c805186",
  1173 => x"da2d86c7",
  1174 => x"2d78802e",
  1175 => x"883880d7",
  1176 => x"ec51a4e9",
  1177 => x"0480d994",
  1178 => x"51afb92d",
  1179 => x"7880dbe0",
  1180 => x"0c02b005",
  1181 => x"0d0402ec",
  1182 => x"050d80dc",
  1183 => x"cc0b80d7",
  1184 => x"e80c80dc",
  1185 => x"cc558075",
  1186 => x"81b72d80",
  1187 => x"d9b80851",
  1188 => x"a2c52dba",
  1189 => x"51a2902d",
  1190 => x"ffb40870",
  1191 => x"8c2a5154",
  1192 => x"8051a2c5",
  1193 => x"2d73902a",
  1194 => x"51a2c52d",
  1195 => x"73882a70",
  1196 => x"81ff0652",
  1197 => x"53a2c52d",
  1198 => x"7381ff06",
  1199 => x"51a2c52d",
  1200 => x"745280dc",
  1201 => x"8851a2f6",
  1202 => x"2d80d7ec",
  1203 => x"51afb92d",
  1204 => x"80d9b808",
  1205 => x"840580d9",
  1206 => x"b80c0294",
  1207 => x"050d0480",
  1208 => x"0b80d9b8",
  1209 => x"0c0402ec",
  1210 => x"050d840b",
  1211 => x"ec0cacf6",
  1212 => x"2da7dc2d",
  1213 => x"81f92d83",
  1214 => x"53acd92d",
  1215 => x"8151858d",
  1216 => x"2dff1353",
  1217 => x"728025f1",
  1218 => x"38840bec",
  1219 => x"0c80d684",
  1220 => x"5186a02d",
  1221 => x"80c1b42d",
  1222 => x"80dbe008",
  1223 => x"802e81a5",
  1224 => x"38a39d51",
  1225 => x"80d4b42d",
  1226 => x"80d69c52",
  1227 => x"80dc8851",
  1228 => x"a2f62d80",
  1229 => x"d7ec51af",
  1230 => x"b92dad98",
  1231 => x"2da8ad2d",
  1232 => x"afcc2d80",
  1233 => x"d8800b80",
  1234 => x"f52d80da",
  1235 => x"9c087081",
  1236 => x"06555654",
  1237 => x"72802e85",
  1238 => x"38738407",
  1239 => x"5474812a",
  1240 => x"70810651",
  1241 => x"5372802e",
  1242 => x"85387382",
  1243 => x"07547482",
  1244 => x"2a708106",
  1245 => x"51537280",
  1246 => x"2e853873",
  1247 => x"81075474",
  1248 => x"832a7081",
  1249 => x"06515372",
  1250 => x"802e8538",
  1251 => x"73880754",
  1252 => x"74842a70",
  1253 => x"81065153",
  1254 => x"72802e85",
  1255 => x"38739007",
  1256 => x"5474852a",
  1257 => x"70810651",
  1258 => x"5372802e",
  1259 => x"853873a0",
  1260 => x"075473fc",
  1261 => x"0c865380",
  1262 => x"dbe00883",
  1263 => x"38845372",
  1264 => x"ec0ca6bd",
  1265 => x"04800b80",
  1266 => x"dbe00c02",
  1267 => x"94050d04",
  1268 => x"71980c04",
  1269 => x"ffb00880",
  1270 => x"dbe00c04",
  1271 => x"810bffb0",
  1272 => x"0c04800b",
  1273 => x"ffb00c04",
  1274 => x"02f8050d",
  1275 => x"ffb40870",
  1276 => x"9fff0651",
  1277 => x"517080da",
  1278 => x"8c082e8c",
  1279 => x"387080da",
  1280 => x"8c0c800b",
  1281 => x"80da880c",
  1282 => x"80da8808",
  1283 => x"51815270",
  1284 => x"87e82e8f",
  1285 => x"387087e8",
  1286 => x"24873871",
  1287 => x"1180da88",
  1288 => x"0c805271",
  1289 => x"80dbe00c",
  1290 => x"0288050d",
  1291 => x"0402e005",
  1292 => x"0da9bb04",
  1293 => x"80dbe008",
  1294 => x"81f02e09",
  1295 => x"81068a38",
  1296 => x"810b80da",
  1297 => x"940ca9bb",
  1298 => x"0480dbe0",
  1299 => x"0881e02e",
  1300 => x"0981068a",
  1301 => x"38810b80",
  1302 => x"da980ca9",
  1303 => x"bb0480db",
  1304 => x"e0085280",
  1305 => x"da980880",
  1306 => x"2e893880",
  1307 => x"dbe00881",
  1308 => x"80055271",
  1309 => x"842c728f",
  1310 => x"06535380",
  1311 => x"da940880",
  1312 => x"2e9a3872",
  1313 => x"842980d9",
  1314 => x"bc057213",
  1315 => x"81712b70",
  1316 => x"09730806",
  1317 => x"730c5153",
  1318 => x"53a9af04",
  1319 => x"72842980",
  1320 => x"d9bc0572",
  1321 => x"1383712b",
  1322 => x"72080772",
  1323 => x"0c535380",
  1324 => x"0b80da98",
  1325 => x"0c800b80",
  1326 => x"da940c80",
  1327 => x"dd9051ab",
  1328 => x"cc2d80db",
  1329 => x"e008ff24",
  1330 => x"feea38a7",
  1331 => x"e82d80db",
  1332 => x"e008802e",
  1333 => x"80ff3881",
  1334 => x"56800b80",
  1335 => x"da900880",
  1336 => x"da8c0880",
  1337 => x"da940857",
  1338 => x"59595577",
  1339 => x"76067777",
  1340 => x"06545271",
  1341 => x"732e80c4",
  1342 => x"387280d9",
  1343 => x"fc1680f5",
  1344 => x"2d70842c",
  1345 => x"718f0652",
  1346 => x"55535473",
  1347 => x"802e9a38",
  1348 => x"72842980",
  1349 => x"d9bc0572",
  1350 => x"1381712b",
  1351 => x"70097308",
  1352 => x"06730c51",
  1353 => x"5353aabc",
  1354 => x"04728429",
  1355 => x"80d9bc05",
  1356 => x"72138371",
  1357 => x"2b720807",
  1358 => x"720c5353",
  1359 => x"75108116",
  1360 => x"56568b75",
  1361 => x"25ffa438",
  1362 => x"7380da94",
  1363 => x"0c80da8c",
  1364 => x"0880da90",
  1365 => x"0c800b80",
  1366 => x"dbe00c02",
  1367 => x"a0050d04",
  1368 => x"02f8050d",
  1369 => x"80d9bc52",
  1370 => x"8f518072",
  1371 => x"70840554",
  1372 => x"0cff1151",
  1373 => x"708025f2",
  1374 => x"38028805",
  1375 => x"0d0402f0",
  1376 => x"050d7551",
  1377 => x"a7e22d70",
  1378 => x"822cfc06",
  1379 => x"80d9bc11",
  1380 => x"72109e06",
  1381 => x"71087072",
  1382 => x"2a708306",
  1383 => x"82742b70",
  1384 => x"09740676",
  1385 => x"0c545156",
  1386 => x"57535153",
  1387 => x"a7dc2d71",
  1388 => x"80dbe00c",
  1389 => x"0290050d",
  1390 => x"0402fc05",
  1391 => x"0d725180",
  1392 => x"710c800b",
  1393 => x"84120c02",
  1394 => x"84050d04",
  1395 => x"02f0050d",
  1396 => x"75700884",
  1397 => x"12085353",
  1398 => x"53ff5471",
  1399 => x"712ea838",
  1400 => x"a7e22d84",
  1401 => x"13087084",
  1402 => x"29148811",
  1403 => x"70087081",
  1404 => x"ff068418",
  1405 => x"08811187",
  1406 => x"06841a0c",
  1407 => x"53515551",
  1408 => x"5151a7dc",
  1409 => x"2d715473",
  1410 => x"80dbe00c",
  1411 => x"0290050d",
  1412 => x"0402f805",
  1413 => x"0da7e22d",
  1414 => x"e008708b",
  1415 => x"2a708106",
  1416 => x"51525270",
  1417 => x"802ea138",
  1418 => x"80dd9008",
  1419 => x"70842980",
  1420 => x"dd980573",
  1421 => x"81ff0671",
  1422 => x"0c515180",
  1423 => x"dd900881",
  1424 => x"11870680",
  1425 => x"dd900c51",
  1426 => x"800b80dd",
  1427 => x"b80ca7d4",
  1428 => x"2da7dc2d",
  1429 => x"0288050d",
  1430 => x"0402fc05",
  1431 => x"0da7e22d",
  1432 => x"810b80dd",
  1433 => x"b80ca7dc",
  1434 => x"2d80ddb8",
  1435 => x"085170f9",
  1436 => x"38028405",
  1437 => x"0d0402fc",
  1438 => x"050d80dd",
  1439 => x"9051abb9",
  1440 => x"2daae02d",
  1441 => x"ac9151a7",
  1442 => x"d02d0284",
  1443 => x"050d0480",
  1444 => x"ddc40880",
  1445 => x"dbe00c04",
  1446 => x"02fc050d",
  1447 => x"810b80da",
  1448 => x"a00c8151",
  1449 => x"858d2d02",
  1450 => x"84050d04",
  1451 => x"02fc050d",
  1452 => x"adb604a8",
  1453 => x"ad2d80f6",
  1454 => x"51aafe2d",
  1455 => x"80dbe008",
  1456 => x"f23880da",
  1457 => x"51aafe2d",
  1458 => x"80dbe008",
  1459 => x"e63880db",
  1460 => x"e00880da",
  1461 => x"a00c80db",
  1462 => x"e0085185",
  1463 => x"8d2d0284",
  1464 => x"050d0402",
  1465 => x"ec050d76",
  1466 => x"54805287",
  1467 => x"0b881580",
  1468 => x"f52d5653",
  1469 => x"74722483",
  1470 => x"38a05372",
  1471 => x"5183842d",
  1472 => x"81128b15",
  1473 => x"80f52d54",
  1474 => x"52727225",
  1475 => x"de380294",
  1476 => x"050d0402",
  1477 => x"f0050d80",
  1478 => x"ddc40854",
  1479 => x"81f92d80",
  1480 => x"0b80ddc8",
  1481 => x"0c730880",
  1482 => x"2e818938",
  1483 => x"820b80db",
  1484 => x"f40c80dd",
  1485 => x"c8088f06",
  1486 => x"80dbf00c",
  1487 => x"73085271",
  1488 => x"832e9638",
  1489 => x"71832689",
  1490 => x"3871812e",
  1491 => x"b038af9d",
  1492 => x"0471852e",
  1493 => x"a038af9d",
  1494 => x"04881480",
  1495 => x"f52d8415",
  1496 => x"0880d6ac",
  1497 => x"53545286",
  1498 => x"a02d7184",
  1499 => x"29137008",
  1500 => x"5252afa1",
  1501 => x"047351ad",
  1502 => x"e32daf9d",
  1503 => x"0480da9c",
  1504 => x"08881508",
  1505 => x"2c708106",
  1506 => x"51527180",
  1507 => x"2e883880",
  1508 => x"d6b051af",
  1509 => x"9a0480d6",
  1510 => x"b45186a0",
  1511 => x"2d841408",
  1512 => x"5186a02d",
  1513 => x"80ddc808",
  1514 => x"810580dd",
  1515 => x"c80c8c14",
  1516 => x"54aea504",
  1517 => x"0290050d",
  1518 => x"047180dd",
  1519 => x"c40cae93",
  1520 => x"2d80ddc8",
  1521 => x"08ff0580",
  1522 => x"ddcc0c04",
  1523 => x"02e8050d",
  1524 => x"80ddc408",
  1525 => x"80ddd008",
  1526 => x"575580f6",
  1527 => x"51aafe2d",
  1528 => x"80dbe008",
  1529 => x"812a7081",
  1530 => x"06515271",
  1531 => x"802ea438",
  1532 => x"aff604a8",
  1533 => x"ad2d80f6",
  1534 => x"51aafe2d",
  1535 => x"80dbe008",
  1536 => x"f23880da",
  1537 => x"a0088132",
  1538 => x"7080daa0",
  1539 => x"0c705252",
  1540 => x"858d2d80",
  1541 => x"0b80ddbc",
  1542 => x"0c800b80",
  1543 => x"ddc00c80",
  1544 => x"daa00883",
  1545 => x"8d3880da",
  1546 => x"51aafe2d",
  1547 => x"80dbe008",
  1548 => x"802e8c38",
  1549 => x"80ddbc08",
  1550 => x"81800780",
  1551 => x"ddbc0c80",
  1552 => x"d951aafe",
  1553 => x"2d80dbe0",
  1554 => x"08802e8c",
  1555 => x"3880ddbc",
  1556 => x"0880c007",
  1557 => x"80ddbc0c",
  1558 => x"819451aa",
  1559 => x"fe2d80db",
  1560 => x"e008802e",
  1561 => x"8b3880dd",
  1562 => x"bc089007",
  1563 => x"80ddbc0c",
  1564 => x"819151aa",
  1565 => x"fe2d80db",
  1566 => x"e008802e",
  1567 => x"8b3880dd",
  1568 => x"bc08a007",
  1569 => x"80ddbc0c",
  1570 => x"81f551aa",
  1571 => x"fe2d80db",
  1572 => x"e008802e",
  1573 => x"8b3880dd",
  1574 => x"bc088107",
  1575 => x"80ddbc0c",
  1576 => x"81f251aa",
  1577 => x"fe2d80db",
  1578 => x"e008802e",
  1579 => x"8b3880dd",
  1580 => x"bc088207",
  1581 => x"80ddbc0c",
  1582 => x"81eb51aa",
  1583 => x"fe2d80db",
  1584 => x"e008802e",
  1585 => x"8b3880dd",
  1586 => x"bc088407",
  1587 => x"80ddbc0c",
  1588 => x"81f451aa",
  1589 => x"fe2d80db",
  1590 => x"e008802e",
  1591 => x"8b3880dd",
  1592 => x"bc088807",
  1593 => x"80ddbc0c",
  1594 => x"80d851aa",
  1595 => x"fe2d80db",
  1596 => x"e008802e",
  1597 => x"8c3880dd",
  1598 => x"c0088180",
  1599 => x"0780ddc0",
  1600 => x"0c9251aa",
  1601 => x"fe2d80db",
  1602 => x"e008802e",
  1603 => x"8c3880dd",
  1604 => x"c00880c0",
  1605 => x"0780ddc0",
  1606 => x"0c9451aa",
  1607 => x"fe2d80db",
  1608 => x"e008802e",
  1609 => x"8b3880dd",
  1610 => x"c0089007",
  1611 => x"80ddc00c",
  1612 => x"9151aafe",
  1613 => x"2d80dbe0",
  1614 => x"08802e8b",
  1615 => x"3880ddc0",
  1616 => x"08a00780",
  1617 => x"ddc00c9d",
  1618 => x"51aafe2d",
  1619 => x"80dbe008",
  1620 => x"802e8b38",
  1621 => x"80ddc008",
  1622 => x"810780dd",
  1623 => x"c00c9b51",
  1624 => x"aafe2d80",
  1625 => x"dbe00880",
  1626 => x"2e8b3880",
  1627 => x"ddc00882",
  1628 => x"0780ddc0",
  1629 => x"0c9c51aa",
  1630 => x"fe2d80db",
  1631 => x"e008802e",
  1632 => x"8b3880dd",
  1633 => x"c0088407",
  1634 => x"80ddc00c",
  1635 => x"a351aafe",
  1636 => x"2d80dbe0",
  1637 => x"08802e8b",
  1638 => x"3880ddc0",
  1639 => x"08880780",
  1640 => x"ddc00c81",
  1641 => x"fd51aafe",
  1642 => x"2d81fa51",
  1643 => x"aafe2db9",
  1644 => x"870481f5",
  1645 => x"51aafe2d",
  1646 => x"80dbe008",
  1647 => x"812a7081",
  1648 => x"06515271",
  1649 => x"802eb338",
  1650 => x"80ddcc08",
  1651 => x"5271802e",
  1652 => x"8a38ff12",
  1653 => x"80ddcc0c",
  1654 => x"b3fa0480",
  1655 => x"ddc80810",
  1656 => x"80ddc808",
  1657 => x"05708429",
  1658 => x"16515288",
  1659 => x"1208802e",
  1660 => x"8938ff51",
  1661 => x"88120852",
  1662 => x"712d81f2",
  1663 => x"51aafe2d",
  1664 => x"80dbe008",
  1665 => x"812a7081",
  1666 => x"06515271",
  1667 => x"802eb438",
  1668 => x"80ddc808",
  1669 => x"ff1180dd",
  1670 => x"cc085653",
  1671 => x"53737225",
  1672 => x"8a388114",
  1673 => x"80ddcc0c",
  1674 => x"b4c30472",
  1675 => x"10137084",
  1676 => x"29165152",
  1677 => x"88120880",
  1678 => x"2e8938fe",
  1679 => x"51881208",
  1680 => x"52712d81",
  1681 => x"fd51aafe",
  1682 => x"2d80dbe0",
  1683 => x"08812a70",
  1684 => x"81065152",
  1685 => x"71802eb1",
  1686 => x"3880ddcc",
  1687 => x"08802e8a",
  1688 => x"38800b80",
  1689 => x"ddcc0cb5",
  1690 => x"890480dd",
  1691 => x"c8081080",
  1692 => x"ddc80805",
  1693 => x"70842916",
  1694 => x"51528812",
  1695 => x"08802e89",
  1696 => x"38fd5188",
  1697 => x"12085271",
  1698 => x"2d81fa51",
  1699 => x"aafe2d80",
  1700 => x"dbe00881",
  1701 => x"2a708106",
  1702 => x"51527180",
  1703 => x"2eb13880",
  1704 => x"ddc808ff",
  1705 => x"11545280",
  1706 => x"ddcc0873",
  1707 => x"25893872",
  1708 => x"80ddcc0c",
  1709 => x"b5cf0471",
  1710 => x"10127084",
  1711 => x"29165152",
  1712 => x"88120880",
  1713 => x"2e8938fc",
  1714 => x"51881208",
  1715 => x"52712d80",
  1716 => x"ddcc0870",
  1717 => x"53547380",
  1718 => x"2e8a388c",
  1719 => x"15ff1555",
  1720 => x"55b5d604",
  1721 => x"820b80db",
  1722 => x"f40c718f",
  1723 => x"0680dbf0",
  1724 => x"0c81eb51",
  1725 => x"aafe2d80",
  1726 => x"dbe00881",
  1727 => x"2a708106",
  1728 => x"51527180",
  1729 => x"2ead3874",
  1730 => x"08852e09",
  1731 => x"8106a438",
  1732 => x"881580f5",
  1733 => x"2dff0552",
  1734 => x"71881681",
  1735 => x"b72d7198",
  1736 => x"2b527180",
  1737 => x"25883880",
  1738 => x"0b881681",
  1739 => x"b72d7451",
  1740 => x"ade32d81",
  1741 => x"f451aafe",
  1742 => x"2d80dbe0",
  1743 => x"08812a70",
  1744 => x"81065152",
  1745 => x"71802eb3",
  1746 => x"38740885",
  1747 => x"2e098106",
  1748 => x"aa388815",
  1749 => x"80f52d81",
  1750 => x"05527188",
  1751 => x"1681b72d",
  1752 => x"7181ff06",
  1753 => x"8b1680f5",
  1754 => x"2d545272",
  1755 => x"72278738",
  1756 => x"72881681",
  1757 => x"b72d7451",
  1758 => x"ade32d80",
  1759 => x"da51aafe",
  1760 => x"2d80dbe0",
  1761 => x"08812a70",
  1762 => x"81065152",
  1763 => x"71802e81",
  1764 => x"ad3880dd",
  1765 => x"c40880dd",
  1766 => x"cc085553",
  1767 => x"73802e8a",
  1768 => x"388c13ff",
  1769 => x"155553b7",
  1770 => x"9c047208",
  1771 => x"5271822e",
  1772 => x"a6387182",
  1773 => x"26893871",
  1774 => x"812eaa38",
  1775 => x"b8be0471",
  1776 => x"832eb438",
  1777 => x"71842e09",
  1778 => x"810680f2",
  1779 => x"38881308",
  1780 => x"51afb92d",
  1781 => x"b8be0480",
  1782 => x"ddcc0851",
  1783 => x"88130852",
  1784 => x"712db8be",
  1785 => x"04810b88",
  1786 => x"14082b80",
  1787 => x"da9c0832",
  1788 => x"80da9c0c",
  1789 => x"b8920488",
  1790 => x"1380f52d",
  1791 => x"81058b14",
  1792 => x"80f52d53",
  1793 => x"54717424",
  1794 => x"83388054",
  1795 => x"73881481",
  1796 => x"b72dae93",
  1797 => x"2db8be04",
  1798 => x"7508802e",
  1799 => x"a4387508",
  1800 => x"51aafe2d",
  1801 => x"80dbe008",
  1802 => x"81065271",
  1803 => x"802e8c38",
  1804 => x"80ddcc08",
  1805 => x"51841608",
  1806 => x"52712d88",
  1807 => x"165675d8",
  1808 => x"38805480",
  1809 => x"0b80dbf4",
  1810 => x"0c738f06",
  1811 => x"80dbf00c",
  1812 => x"a0527380",
  1813 => x"ddcc082e",
  1814 => x"09810699",
  1815 => x"3880ddc8",
  1816 => x"08ff0574",
  1817 => x"32700981",
  1818 => x"05707207",
  1819 => x"9f2a9171",
  1820 => x"31515153",
  1821 => x"53715183",
  1822 => x"842d8114",
  1823 => x"548e7425",
  1824 => x"c23880da",
  1825 => x"a0085271",
  1826 => x"80dbe00c",
  1827 => x"0298050d",
  1828 => x"0402f405",
  1829 => x"0dd45281",
  1830 => x"ff720c71",
  1831 => x"085381ff",
  1832 => x"720c7288",
  1833 => x"2b83fe80",
  1834 => x"06720870",
  1835 => x"81ff0651",
  1836 => x"525381ff",
  1837 => x"720c7271",
  1838 => x"07882b72",
  1839 => x"087081ff",
  1840 => x"06515253",
  1841 => x"81ff720c",
  1842 => x"72710788",
  1843 => x"2b720870",
  1844 => x"81ff0672",
  1845 => x"0780dbe0",
  1846 => x"0c525302",
  1847 => x"8c050d04",
  1848 => x"02f4050d",
  1849 => x"74767181",
  1850 => x"ff06d40c",
  1851 => x"535380dd",
  1852 => x"d4088538",
  1853 => x"71892b52",
  1854 => x"71982ad4",
  1855 => x"0c71902a",
  1856 => x"7081ff06",
  1857 => x"d40c5171",
  1858 => x"882a7081",
  1859 => x"ff06d40c",
  1860 => x"517181ff",
  1861 => x"06d40c72",
  1862 => x"902a7081",
  1863 => x"ff06d40c",
  1864 => x"51d40870",
  1865 => x"81ff0651",
  1866 => x"5182b8bf",
  1867 => x"527081ff",
  1868 => x"2e098106",
  1869 => x"943881ff",
  1870 => x"0bd40cd4",
  1871 => x"087081ff",
  1872 => x"06ff1454",
  1873 => x"515171e5",
  1874 => x"387080db",
  1875 => x"e00c028c",
  1876 => x"050d0402",
  1877 => x"fc050d81",
  1878 => x"c75181ff",
  1879 => x"0bd40cff",
  1880 => x"11517080",
  1881 => x"25f43802",
  1882 => x"84050d04",
  1883 => x"02f4050d",
  1884 => x"81ff0bd4",
  1885 => x"0c935380",
  1886 => x"5287fc80",
  1887 => x"c151b9e0",
  1888 => x"2d80dbe0",
  1889 => x"088b3881",
  1890 => x"ff0bd40c",
  1891 => x"8153bb9a",
  1892 => x"04bad32d",
  1893 => x"ff135372",
  1894 => x"de387280",
  1895 => x"dbe00c02",
  1896 => x"8c050d04",
  1897 => x"02ec050d",
  1898 => x"810b80dd",
  1899 => x"d40c8454",
  1900 => x"d008708f",
  1901 => x"2a708106",
  1902 => x"51515372",
  1903 => x"f33872d0",
  1904 => x"0cbad32d",
  1905 => x"80d6b851",
  1906 => x"86a02dd0",
  1907 => x"08708f2a",
  1908 => x"70810651",
  1909 => x"515372f3",
  1910 => x"38810bd0",
  1911 => x"0cb15380",
  1912 => x"5284d480",
  1913 => x"c051b9e0",
  1914 => x"2d80dbe0",
  1915 => x"08812e93",
  1916 => x"3872822e",
  1917 => x"bf38ff13",
  1918 => x"5372e438",
  1919 => x"ff145473",
  1920 => x"ffae38ba",
  1921 => x"d32d83aa",
  1922 => x"52849c80",
  1923 => x"c851b9e0",
  1924 => x"2d80dbe0",
  1925 => x"08812e09",
  1926 => x"81069338",
  1927 => x"b9912d80",
  1928 => x"dbe00883",
  1929 => x"ffff0653",
  1930 => x"7283aa2e",
  1931 => x"9f38baec",
  1932 => x"2dbcc704",
  1933 => x"80d6c451",
  1934 => x"86a02d80",
  1935 => x"53be9c04",
  1936 => x"80d6dc51",
  1937 => x"86a02d80",
  1938 => x"54bded04",
  1939 => x"81ff0bd4",
  1940 => x"0cb154ba",
  1941 => x"d32d8fcf",
  1942 => x"53805287",
  1943 => x"fc80f751",
  1944 => x"b9e02d80",
  1945 => x"dbe00855",
  1946 => x"80dbe008",
  1947 => x"812e0981",
  1948 => x"069c3881",
  1949 => x"ff0bd40c",
  1950 => x"820a5284",
  1951 => x"9c80e951",
  1952 => x"b9e02d80",
  1953 => x"dbe00880",
  1954 => x"2e8d38ba",
  1955 => x"d32dff13",
  1956 => x"5372c638",
  1957 => x"bde00481",
  1958 => x"ff0bd40c",
  1959 => x"80dbe008",
  1960 => x"5287fc80",
  1961 => x"fa51b9e0",
  1962 => x"2d80dbe0",
  1963 => x"08b23881",
  1964 => x"ff0bd40c",
  1965 => x"d4085381",
  1966 => x"ff0bd40c",
  1967 => x"81ff0bd4",
  1968 => x"0c81ff0b",
  1969 => x"d40c81ff",
  1970 => x"0bd40c72",
  1971 => x"862a7081",
  1972 => x"06765651",
  1973 => x"53729638",
  1974 => x"80dbe008",
  1975 => x"54bded04",
  1976 => x"73822efe",
  1977 => x"db38ff14",
  1978 => x"5473fee7",
  1979 => x"387380dd",
  1980 => x"d40c738b",
  1981 => x"38815287",
  1982 => x"fc80d051",
  1983 => x"b9e02d81",
  1984 => x"ff0bd40c",
  1985 => x"d008708f",
  1986 => x"2a708106",
  1987 => x"51515372",
  1988 => x"f33872d0",
  1989 => x"0c81ff0b",
  1990 => x"d40c8153",
  1991 => x"7280dbe0",
  1992 => x"0c029405",
  1993 => x"0d0402e8",
  1994 => x"050d7855",
  1995 => x"805681ff",
  1996 => x"0bd40cd0",
  1997 => x"08708f2a",
  1998 => x"70810651",
  1999 => x"515372f3",
  2000 => x"3882810b",
  2001 => x"d00c81ff",
  2002 => x"0bd40c77",
  2003 => x"5287fc80",
  2004 => x"d151b9e0",
  2005 => x"2d80dbc6",
  2006 => x"df5480db",
  2007 => x"e008802e",
  2008 => x"8b3880d6",
  2009 => x"fc5186a0",
  2010 => x"2dbfc004",
  2011 => x"81ff0bd4",
  2012 => x"0cd40870",
  2013 => x"81ff0651",
  2014 => x"537281fe",
  2015 => x"2e098106",
  2016 => x"9e3880ff",
  2017 => x"53b9912d",
  2018 => x"80dbe008",
  2019 => x"75708405",
  2020 => x"570cff13",
  2021 => x"53728025",
  2022 => x"ec388156",
  2023 => x"bfa504ff",
  2024 => x"145473c8",
  2025 => x"3881ff0b",
  2026 => x"d40c81ff",
  2027 => x"0bd40cd0",
  2028 => x"08708f2a",
  2029 => x"70810651",
  2030 => x"515372f3",
  2031 => x"3872d00c",
  2032 => x"7580dbe0",
  2033 => x"0c029805",
  2034 => x"0d0402e8",
  2035 => x"050d7779",
  2036 => x"7b585555",
  2037 => x"80537276",
  2038 => x"25a43874",
  2039 => x"70810556",
  2040 => x"80f52d74",
  2041 => x"70810556",
  2042 => x"80f52d52",
  2043 => x"5271712e",
  2044 => x"87388151",
  2045 => x"80c08004",
  2046 => x"811353bf",
  2047 => x"d6048051",
  2048 => x"7080dbe0",
  2049 => x"0c029805",
  2050 => x"0d0402ec",
  2051 => x"050d7655",
  2052 => x"74802e80",
  2053 => x"c4389a15",
  2054 => x"80e02d51",
  2055 => x"80ceb82d",
  2056 => x"80dbe008",
  2057 => x"80dbe008",
  2058 => x"80e4880c",
  2059 => x"80dbe008",
  2060 => x"545480e3",
  2061 => x"e408802e",
  2062 => x"9b389415",
  2063 => x"80e02d51",
  2064 => x"80ceb82d",
  2065 => x"80dbe008",
  2066 => x"902b83ff",
  2067 => x"f00a0670",
  2068 => x"75075153",
  2069 => x"7280e488",
  2070 => x"0c80e488",
  2071 => x"08537280",
  2072 => x"2e9e3880",
  2073 => x"e3dc08fe",
  2074 => x"14712980",
  2075 => x"e3f00805",
  2076 => x"80e48c0c",
  2077 => x"70842b80",
  2078 => x"e3e80c54",
  2079 => x"80c1af04",
  2080 => x"80e3f408",
  2081 => x"80e4880c",
  2082 => x"80e3f808",
  2083 => x"80e48c0c",
  2084 => x"80e3e408",
  2085 => x"802e8c38",
  2086 => x"80e3dc08",
  2087 => x"842b5380",
  2088 => x"c1aa0480",
  2089 => x"e3fc0884",
  2090 => x"2b537280",
  2091 => x"e3e80c02",
  2092 => x"94050d04",
  2093 => x"02d8050d",
  2094 => x"800b80e3",
  2095 => x"e40c8454",
  2096 => x"bba42d80",
  2097 => x"dbe00880",
  2098 => x"2e983880",
  2099 => x"ddd85280",
  2100 => x"51bea62d",
  2101 => x"80dbe008",
  2102 => x"802e8738",
  2103 => x"fe5480c1",
  2104 => x"ea04ff14",
  2105 => x"54738024",
  2106 => x"d738738e",
  2107 => x"3880d78c",
  2108 => x"5186a02d",
  2109 => x"735580c7",
  2110 => x"c8048056",
  2111 => x"810b80e4",
  2112 => x"900c8853",
  2113 => x"80d7a052",
  2114 => x"80de8e51",
  2115 => x"bfca2d80",
  2116 => x"dbe00876",
  2117 => x"2e098106",
  2118 => x"893880db",
  2119 => x"e00880e4",
  2120 => x"900c8853",
  2121 => x"80d7ac52",
  2122 => x"80deaa51",
  2123 => x"bfca2d80",
  2124 => x"dbe00889",
  2125 => x"3880dbe0",
  2126 => x"0880e490",
  2127 => x"0c80e490",
  2128 => x"08802e81",
  2129 => x"843880e1",
  2130 => x"9e0b80f5",
  2131 => x"2d80e19f",
  2132 => x"0b80f52d",
  2133 => x"71982b71",
  2134 => x"902b0780",
  2135 => x"e1a00b80",
  2136 => x"f52d7088",
  2137 => x"2b720780",
  2138 => x"e1a10b80",
  2139 => x"f52d7107",
  2140 => x"80e1d60b",
  2141 => x"80f52d80",
  2142 => x"e1d70b80",
  2143 => x"f52d7188",
  2144 => x"2b07535f",
  2145 => x"54525a56",
  2146 => x"57557381",
  2147 => x"abaa2e09",
  2148 => x"81069038",
  2149 => x"755180ce",
  2150 => x"872d80db",
  2151 => x"e0085680",
  2152 => x"c3b20473",
  2153 => x"82d4d52e",
  2154 => x"893880d7",
  2155 => x"b85180c3",
  2156 => x"ff0480dd",
  2157 => x"d8527551",
  2158 => x"bea62d80",
  2159 => x"dbe00855",
  2160 => x"80dbe008",
  2161 => x"802e8480",
  2162 => x"38885380",
  2163 => x"d7ac5280",
  2164 => x"deaa51bf",
  2165 => x"ca2d80db",
  2166 => x"e0088b38",
  2167 => x"810b80e3",
  2168 => x"e40c80c4",
  2169 => x"86048853",
  2170 => x"80d7a052",
  2171 => x"80de8e51",
  2172 => x"bfca2d80",
  2173 => x"dbe00880",
  2174 => x"2e8c3880",
  2175 => x"d7cc5186",
  2176 => x"a02d80c4",
  2177 => x"e50480e1",
  2178 => x"d60b80f5",
  2179 => x"2d547380",
  2180 => x"d52e0981",
  2181 => x"0680ce38",
  2182 => x"80e1d70b",
  2183 => x"80f52d54",
  2184 => x"7381aa2e",
  2185 => x"098106bd",
  2186 => x"38800b80",
  2187 => x"ddd80b80",
  2188 => x"f52d5654",
  2189 => x"7481e92e",
  2190 => x"83388154",
  2191 => x"7481eb2e",
  2192 => x"8c388055",
  2193 => x"73752e09",
  2194 => x"810682fc",
  2195 => x"3880dde3",
  2196 => x"0b80f52d",
  2197 => x"55748e38",
  2198 => x"80dde40b",
  2199 => x"80f52d54",
  2200 => x"73822e87",
  2201 => x"38805580",
  2202 => x"c7c80480",
  2203 => x"dde50b80",
  2204 => x"f52d7080",
  2205 => x"e3dc0cff",
  2206 => x"0580e3e0",
  2207 => x"0c80dde6",
  2208 => x"0b80f52d",
  2209 => x"80dde70b",
  2210 => x"80f52d58",
  2211 => x"76057782",
  2212 => x"80290570",
  2213 => x"80e3ec0c",
  2214 => x"80dde80b",
  2215 => x"80f52d70",
  2216 => x"80e4800c",
  2217 => x"80e3e408",
  2218 => x"59575876",
  2219 => x"802e81b8",
  2220 => x"38885380",
  2221 => x"d7ac5280",
  2222 => x"deaa51bf",
  2223 => x"ca2d80db",
  2224 => x"e0088284",
  2225 => x"3880e3dc",
  2226 => x"0870842b",
  2227 => x"80e3e80c",
  2228 => x"7080e3fc",
  2229 => x"0c80ddfd",
  2230 => x"0b80f52d",
  2231 => x"80ddfc0b",
  2232 => x"80f52d71",
  2233 => x"82802905",
  2234 => x"80ddfe0b",
  2235 => x"80f52d70",
  2236 => x"84808029",
  2237 => x"1280ddff",
  2238 => x"0b80f52d",
  2239 => x"7081800a",
  2240 => x"29127080",
  2241 => x"e4840c80",
  2242 => x"e4800871",
  2243 => x"2980e3ec",
  2244 => x"08057080",
  2245 => x"e3f00c80",
  2246 => x"de850b80",
  2247 => x"f52d80de",
  2248 => x"840b80f5",
  2249 => x"2d718280",
  2250 => x"290580de",
  2251 => x"860b80f5",
  2252 => x"2d708480",
  2253 => x"80291280",
  2254 => x"de870b80",
  2255 => x"f52d7098",
  2256 => x"2b81f00a",
  2257 => x"06720570",
  2258 => x"80e3f40c",
  2259 => x"fe117e29",
  2260 => x"770580e3",
  2261 => x"f80c5259",
  2262 => x"5243545e",
  2263 => x"51525952",
  2264 => x"5d575957",
  2265 => x"80c7c004",
  2266 => x"80ddea0b",
  2267 => x"80f52d80",
  2268 => x"dde90b80",
  2269 => x"f52d7182",
  2270 => x"80290570",
  2271 => x"80e3e80c",
  2272 => x"70a02983",
  2273 => x"ff057089",
  2274 => x"2a7080e3",
  2275 => x"fc0c80dd",
  2276 => x"ef0b80f5",
  2277 => x"2d80ddee",
  2278 => x"0b80f52d",
  2279 => x"71828029",
  2280 => x"057080e4",
  2281 => x"840c7b71",
  2282 => x"291e7080",
  2283 => x"e3f80c7d",
  2284 => x"80e3f40c",
  2285 => x"730580e3",
  2286 => x"f00c555e",
  2287 => x"51515555",
  2288 => x"805180c0",
  2289 => x"8a2d8155",
  2290 => x"7480dbe0",
  2291 => x"0c02a805",
  2292 => x"0d0402ec",
  2293 => x"050d7670",
  2294 => x"872c7180",
  2295 => x"ff065556",
  2296 => x"5480e3e4",
  2297 => x"088a3873",
  2298 => x"882c7481",
  2299 => x"ff065455",
  2300 => x"80ddd852",
  2301 => x"80e3ec08",
  2302 => x"1551bea6",
  2303 => x"2d80dbe0",
  2304 => x"085480db",
  2305 => x"e008802e",
  2306 => x"bb3880e3",
  2307 => x"e408802e",
  2308 => x"9c387284",
  2309 => x"2980ddd8",
  2310 => x"05700852",
  2311 => x"5380ce87",
  2312 => x"2d80dbe0",
  2313 => x"08f00a06",
  2314 => x"5380c8c2",
  2315 => x"04721080",
  2316 => x"ddd80570",
  2317 => x"80e02d52",
  2318 => x"5380ceb8",
  2319 => x"2d80dbe0",
  2320 => x"08537254",
  2321 => x"7380dbe0",
  2322 => x"0c029405",
  2323 => x"0d0402e0",
  2324 => x"050d7970",
  2325 => x"842c80e4",
  2326 => x"8c080571",
  2327 => x"8f065255",
  2328 => x"53728a38",
  2329 => x"80ddd852",
  2330 => x"7351bea6",
  2331 => x"2d72a029",
  2332 => x"80ddd805",
  2333 => x"54807480",
  2334 => x"f52d5653",
  2335 => x"74732e83",
  2336 => x"38815374",
  2337 => x"81e52e81",
  2338 => x"f5388170",
  2339 => x"74065458",
  2340 => x"72802e81",
  2341 => x"e9388b14",
  2342 => x"80f52d70",
  2343 => x"832a7906",
  2344 => x"5856769c",
  2345 => x"3880daa4",
  2346 => x"08537289",
  2347 => x"387280e1",
  2348 => x"d80b81b7",
  2349 => x"2d7680da",
  2350 => x"a40c7353",
  2351 => x"80cb8004",
  2352 => x"758f2e09",
  2353 => x"810681b6",
  2354 => x"38749f06",
  2355 => x"8d2980e1",
  2356 => x"cb115153",
  2357 => x"811480f5",
  2358 => x"2d737081",
  2359 => x"055581b7",
  2360 => x"2d831480",
  2361 => x"f52d7370",
  2362 => x"81055581",
  2363 => x"b72d8514",
  2364 => x"80f52d73",
  2365 => x"70810555",
  2366 => x"81b72d87",
  2367 => x"1480f52d",
  2368 => x"73708105",
  2369 => x"5581b72d",
  2370 => x"891480f5",
  2371 => x"2d737081",
  2372 => x"055581b7",
  2373 => x"2d8e1480",
  2374 => x"f52d7370",
  2375 => x"81055581",
  2376 => x"b72d9014",
  2377 => x"80f52d73",
  2378 => x"70810555",
  2379 => x"81b72d92",
  2380 => x"1480f52d",
  2381 => x"73708105",
  2382 => x"5581b72d",
  2383 => x"941480f5",
  2384 => x"2d737081",
  2385 => x"055581b7",
  2386 => x"2d961480",
  2387 => x"f52d7370",
  2388 => x"81055581",
  2389 => x"b72d9814",
  2390 => x"80f52d73",
  2391 => x"70810555",
  2392 => x"81b72d9c",
  2393 => x"1480f52d",
  2394 => x"73708105",
  2395 => x"5581b72d",
  2396 => x"9e1480f5",
  2397 => x"2d7381b7",
  2398 => x"2d7780da",
  2399 => x"a40c8053",
  2400 => x"7280dbe0",
  2401 => x"0c02a005",
  2402 => x"0d0402cc",
  2403 => x"050d7e60",
  2404 => x"5e5a800b",
  2405 => x"80e48808",
  2406 => x"80e48c08",
  2407 => x"595c5680",
  2408 => x"5880e3e8",
  2409 => x"08782e81",
  2410 => x"bc38778f",
  2411 => x"06a01757",
  2412 => x"54739138",
  2413 => x"80ddd852",
  2414 => x"76518117",
  2415 => x"57bea62d",
  2416 => x"80ddd856",
  2417 => x"807680f5",
  2418 => x"2d565474",
  2419 => x"742e8338",
  2420 => x"81547481",
  2421 => x"e52e8181",
  2422 => x"38817075",
  2423 => x"06555c73",
  2424 => x"802e80f5",
  2425 => x"388b1680",
  2426 => x"f52d9806",
  2427 => x"597880e9",
  2428 => x"388b537c",
  2429 => x"527551bf",
  2430 => x"ca2d80db",
  2431 => x"e00880d9",
  2432 => x"389c1608",
  2433 => x"5180ce87",
  2434 => x"2d80dbe0",
  2435 => x"08841b0c",
  2436 => x"9a1680e0",
  2437 => x"2d5180ce",
  2438 => x"b82d80db",
  2439 => x"e00880db",
  2440 => x"e008881c",
  2441 => x"0c80dbe0",
  2442 => x"08555580",
  2443 => x"e3e40880",
  2444 => x"2e9a3894",
  2445 => x"1680e02d",
  2446 => x"5180ceb8",
  2447 => x"2d80dbe0",
  2448 => x"08902b83",
  2449 => x"fff00a06",
  2450 => x"70165154",
  2451 => x"73881b0c",
  2452 => x"787a0c7b",
  2453 => x"5480cda3",
  2454 => x"04811858",
  2455 => x"80e3e808",
  2456 => x"7826fec6",
  2457 => x"3880e3e4",
  2458 => x"08802eb5",
  2459 => x"387a5180",
  2460 => x"c7d22d80",
  2461 => x"dbe00880",
  2462 => x"dbe00880",
  2463 => x"fffffff8",
  2464 => x"06555b73",
  2465 => x"80ffffff",
  2466 => x"f82e9638",
  2467 => x"80dbe008",
  2468 => x"fe0580e3",
  2469 => x"dc082980",
  2470 => x"e3f00805",
  2471 => x"5780cb9f",
  2472 => x"04805473",
  2473 => x"80dbe00c",
  2474 => x"02b4050d",
  2475 => x"0402f405",
  2476 => x"0d747008",
  2477 => x"8105710c",
  2478 => x"700880e3",
  2479 => x"e0080653",
  2480 => x"53719038",
  2481 => x"88130851",
  2482 => x"80c7d22d",
  2483 => x"80dbe008",
  2484 => x"88140c81",
  2485 => x"0b80dbe0",
  2486 => x"0c028c05",
  2487 => x"0d0402f0",
  2488 => x"050d7588",
  2489 => x"1108fe05",
  2490 => x"80e3dc08",
  2491 => x"2980e3f0",
  2492 => x"08117208",
  2493 => x"80e3e008",
  2494 => x"06057955",
  2495 => x"535454be",
  2496 => x"a62d0290",
  2497 => x"050d0402",
  2498 => x"f4050d74",
  2499 => x"70882a83",
  2500 => x"fe800670",
  2501 => x"72982a07",
  2502 => x"72882b87",
  2503 => x"fc808006",
  2504 => x"73982b81",
  2505 => x"f00a0671",
  2506 => x"73070780",
  2507 => x"dbe00c56",
  2508 => x"51535102",
  2509 => x"8c050d04",
  2510 => x"02f8050d",
  2511 => x"028e0580",
  2512 => x"f52d7488",
  2513 => x"2b077083",
  2514 => x"ffff0680",
  2515 => x"dbe00c51",
  2516 => x"0288050d",
  2517 => x"0402f405",
  2518 => x"0d747678",
  2519 => x"53545280",
  2520 => x"71259738",
  2521 => x"72708105",
  2522 => x"5480f52d",
  2523 => x"72708105",
  2524 => x"5481b72d",
  2525 => x"ff115170",
  2526 => x"eb388072",
  2527 => x"81b72d02",
  2528 => x"8c050d04",
  2529 => x"02e8050d",
  2530 => x"77568070",
  2531 => x"56547376",
  2532 => x"24b73880",
  2533 => x"e3e80874",
  2534 => x"2eaf3873",
  2535 => x"5180c8ce",
  2536 => x"2d80dbe0",
  2537 => x"0880dbe0",
  2538 => x"08098105",
  2539 => x"7080dbe0",
  2540 => x"08079f2a",
  2541 => x"77058117",
  2542 => x"57575353",
  2543 => x"74762489",
  2544 => x"3880e3e8",
  2545 => x"087426d3",
  2546 => x"387280db",
  2547 => x"e00c0298",
  2548 => x"050d0402",
  2549 => x"f0050d80",
  2550 => x"dbdc0816",
  2551 => x"5180cf84",
  2552 => x"2d80dbe0",
  2553 => x"08802ea0",
  2554 => x"388b5380",
  2555 => x"dbe00852",
  2556 => x"80e1d851",
  2557 => x"80ced52d",
  2558 => x"80e49408",
  2559 => x"5473802e",
  2560 => x"873880e1",
  2561 => x"d851732d",
  2562 => x"0290050d",
  2563 => x"0402dc05",
  2564 => x"0d80705a",
  2565 => x"557480db",
  2566 => x"dc0825b5",
  2567 => x"3880e3e8",
  2568 => x"08752ead",
  2569 => x"38785180",
  2570 => x"c8ce2d80",
  2571 => x"dbe00809",
  2572 => x"81057080",
  2573 => x"dbe00807",
  2574 => x"9f2a7605",
  2575 => x"811b5b56",
  2576 => x"547480db",
  2577 => x"dc082589",
  2578 => x"3880e3e8",
  2579 => x"087926d5",
  2580 => x"38805578",
  2581 => x"80e3e808",
  2582 => x"2781e438",
  2583 => x"785180c8",
  2584 => x"ce2d80db",
  2585 => x"e008802e",
  2586 => x"81b43880",
  2587 => x"dbe0088b",
  2588 => x"0580f52d",
  2589 => x"70842a70",
  2590 => x"81067710",
  2591 => x"78842b80",
  2592 => x"e1d80b80",
  2593 => x"f52d5c5c",
  2594 => x"53515556",
  2595 => x"73802e80",
  2596 => x"ce387416",
  2597 => x"822b80d2",
  2598 => x"e30b80da",
  2599 => x"b0120c54",
  2600 => x"77753110",
  2601 => x"80e49811",
  2602 => x"55569074",
  2603 => x"70810556",
  2604 => x"81b72da0",
  2605 => x"7481b72d",
  2606 => x"7681ff06",
  2607 => x"81165854",
  2608 => x"73802e8b",
  2609 => x"389c5380",
  2610 => x"e1d85280",
  2611 => x"d1d6048b",
  2612 => x"5380dbe0",
  2613 => x"085280e4",
  2614 => x"9a165180",
  2615 => x"d2940474",
  2616 => x"16822b80",
  2617 => x"cfd30b80",
  2618 => x"dab0120c",
  2619 => x"547681ff",
  2620 => x"06811658",
  2621 => x"5473802e",
  2622 => x"8b389c53",
  2623 => x"80e1d852",
  2624 => x"80d28b04",
  2625 => x"8b5380db",
  2626 => x"e0085277",
  2627 => x"75311080",
  2628 => x"e4980551",
  2629 => x"765580ce",
  2630 => x"d52d80d2",
  2631 => x"b3047490",
  2632 => x"29753170",
  2633 => x"1080e498",
  2634 => x"05515480",
  2635 => x"dbe00874",
  2636 => x"81b72d81",
  2637 => x"1959748b",
  2638 => x"24a43880",
  2639 => x"d0d30474",
  2640 => x"90297531",
  2641 => x"701080e4",
  2642 => x"98058c77",
  2643 => x"31575154",
  2644 => x"807481b7",
  2645 => x"2d9e14ff",
  2646 => x"16565474",
  2647 => x"f33802a4",
  2648 => x"050d0402",
  2649 => x"fc050d80",
  2650 => x"dbdc0813",
  2651 => x"5180cf84",
  2652 => x"2d80dbe0",
  2653 => x"08802e8a",
  2654 => x"3880dbe0",
  2655 => x"085180c0",
  2656 => x"8a2d800b",
  2657 => x"80dbdc0c",
  2658 => x"80d08d2d",
  2659 => x"ae932d02",
  2660 => x"84050d04",
  2661 => x"02fc050d",
  2662 => x"725170fd",
  2663 => x"2eb23870",
  2664 => x"fd248b38",
  2665 => x"70fc2e80",
  2666 => x"d03880d4",
  2667 => x"830470fe",
  2668 => x"2eb93870",
  2669 => x"ff2e0981",
  2670 => x"0680c838",
  2671 => x"80dbdc08",
  2672 => x"5170802e",
  2673 => x"be38ff11",
  2674 => x"80dbdc0c",
  2675 => x"80d48304",
  2676 => x"80dbdc08",
  2677 => x"f0057080",
  2678 => x"dbdc0c51",
  2679 => x"708025a3",
  2680 => x"38800b80",
  2681 => x"dbdc0c80",
  2682 => x"d4830480",
  2683 => x"dbdc0881",
  2684 => x"0580dbdc",
  2685 => x"0c80d483",
  2686 => x"0480dbdc",
  2687 => x"08900580",
  2688 => x"dbdc0c80",
  2689 => x"d08d2dae",
  2690 => x"932d0284",
  2691 => x"050d0402",
  2692 => x"fc050d80",
  2693 => x"0b80dbdc",
  2694 => x"0c80d08d",
  2695 => x"2dad8f2d",
  2696 => x"80dbe008",
  2697 => x"80dbcc0c",
  2698 => x"80daa851",
  2699 => x"afb92d02",
  2700 => x"84050d04",
  2701 => x"7180e494",
  2702 => x"0c040000",
  2703 => x"00ffffff",
  2704 => x"ff00ffff",
  2705 => x"ffff00ff",
  2706 => x"ffffff00",
  2707 => x"30313233",
  2708 => x"34353637",
  2709 => x"38394142",
  2710 => x"43444546",
  2711 => x"00000000",
  2712 => x"44656275",
  2713 => x"67000000",
  2714 => x"52657365",
  2715 => x"74000000",
  2716 => x"5363616e",
  2717 => x"6c696e65",
  2718 => x"73000000",
  2719 => x"50414c20",
  2720 => x"2f204e54",
  2721 => x"53430000",
  2722 => x"436f6c6f",
  2723 => x"72000000",
  2724 => x"44696666",
  2725 => x"6963756c",
  2726 => x"74792041",
  2727 => x"00000000",
  2728 => x"44696666",
  2729 => x"6963756c",
  2730 => x"74792042",
  2731 => x"00000000",
  2732 => x"53757065",
  2733 => x"72636869",
  2734 => x"7020696e",
  2735 => x"20636172",
  2736 => x"74726964",
  2737 => x"67650000",
  2738 => x"53656c65",
  2739 => x"63740000",
  2740 => x"53746172",
  2741 => x"74000000",
  2742 => x"4c6f6164",
  2743 => x"20524f4d",
  2744 => x"20100000",
  2745 => x"45786974",
  2746 => x"00000000",
  2747 => x"524f4d20",
  2748 => x"6c6f6164",
  2749 => x"696e6720",
  2750 => x"6661696c",
  2751 => x"65640000",
  2752 => x"4f4b0000",
  2753 => x"496e6974",
  2754 => x"69616c69",
  2755 => x"7a696e67",
  2756 => x"20534420",
  2757 => x"63617264",
  2758 => x"0a000000",
  2759 => x"436f6c6c",
  2760 => x"6563746f",
  2761 => x"72566973",
  2762 => x"696f6e00",
  2763 => x"16200000",
  2764 => x"14200000",
  2765 => x"15200000",
  2766 => x"53442069",
  2767 => x"6e69742e",
  2768 => x"2e2e0a00",
  2769 => x"53442063",
  2770 => x"61726420",
  2771 => x"72657365",
  2772 => x"74206661",
  2773 => x"696c6564",
  2774 => x"210a0000",
  2775 => x"53444843",
  2776 => x"20657272",
  2777 => x"6f72210a",
  2778 => x"00000000",
  2779 => x"57726974",
  2780 => x"65206661",
  2781 => x"696c6564",
  2782 => x"0a000000",
  2783 => x"52656164",
  2784 => x"20666169",
  2785 => x"6c65640a",
  2786 => x"00000000",
  2787 => x"43617264",
  2788 => x"20696e69",
  2789 => x"74206661",
  2790 => x"696c6564",
  2791 => x"0a000000",
  2792 => x"46415431",
  2793 => x"36202020",
  2794 => x"00000000",
  2795 => x"46415433",
  2796 => x"32202020",
  2797 => x"00000000",
  2798 => x"4e6f2070",
  2799 => x"61727469",
  2800 => x"74696f6e",
  2801 => x"20736967",
  2802 => x"0a000000",
  2803 => x"42616420",
  2804 => x"70617274",
  2805 => x"0a000000",
  2806 => x"4261636b",
  2807 => x"00000000",
  2808 => x"00000002",
  2809 => x"00002a4c",
  2810 => x"00002e4c",
  2811 => x"00000002",
  2812 => x"00002e08",
  2813 => x"000012df",
  2814 => x"00000002",
  2815 => x"00002a60",
  2816 => x"00001276",
  2817 => x"00000002",
  2818 => x"00002a68",
  2819 => x"0000035a",
  2820 => x"00000001",
  2821 => x"00002a70",
  2822 => x"00000000",
  2823 => x"00000001",
  2824 => x"00002a7c",
  2825 => x"00000001",
  2826 => x"00000001",
  2827 => x"00002a88",
  2828 => x"00000002",
  2829 => x"00000001",
  2830 => x"00002a90",
  2831 => x"00000003",
  2832 => x"00000001",
  2833 => x"00002aa0",
  2834 => x"00000004",
  2835 => x"00000001",
  2836 => x"00002ab0",
  2837 => x"00000005",
  2838 => x"00000002",
  2839 => x"00002ac8",
  2840 => x"0000036e",
  2841 => x"00000002",
  2842 => x"00002ad0",
  2843 => x"00000a3f",
  2844 => x"00000002",
  2845 => x"00002ad8",
  2846 => x"00002a0f",
  2847 => x"00000002",
  2848 => x"00002ae4",
  2849 => x"000016ac",
  2850 => x"00000000",
  2851 => x"00000000",
  2852 => x"00000000",
  2853 => x"00000004",
  2854 => x"00002aec",
  2855 => x"00002c94",
  2856 => x"00000004",
  2857 => x"00002b00",
  2858 => x"00002bec",
  2859 => x"00000000",
  2860 => x"00000000",
  2861 => x"00000000",
  2862 => x"00000000",
  2863 => x"00000000",
  2864 => x"00000000",
  2865 => x"00000000",
  2866 => x"00000000",
  2867 => x"00000000",
  2868 => x"00000000",
  2869 => x"00000000",
  2870 => x"00000000",
  2871 => x"00000000",
  2872 => x"00000000",
  2873 => x"00000000",
  2874 => x"00000000",
  2875 => x"00000000",
  2876 => x"00000000",
  2877 => x"00000000",
  2878 => x"00000000",
  2879 => x"76f55a1c",
  2880 => x"f21c1c1c",
  2881 => x"1c1c1c1c",
  2882 => x"00000000",
  2883 => x"00000fff",
  2884 => x"00000fff",
  2885 => x"00000000",
  2886 => x"00000000",
  2887 => x"00000006",
  2888 => x"00000000",
  2889 => x"00000000",
  2890 => x"00000002",
  2891 => x"00003218",
  2892 => x"000027d3",
  2893 => x"00000002",
  2894 => x"00003236",
  2895 => x"000027d3",
  2896 => x"00000002",
  2897 => x"00003254",
  2898 => x"000027d3",
  2899 => x"00000002",
  2900 => x"00003272",
  2901 => x"000027d3",
  2902 => x"00000002",
  2903 => x"00003290",
  2904 => x"000027d3",
  2905 => x"00000002",
  2906 => x"000032ae",
  2907 => x"000027d3",
  2908 => x"00000002",
  2909 => x"000032cc",
  2910 => x"000027d3",
  2911 => x"00000002",
  2912 => x"000032ea",
  2913 => x"000027d3",
  2914 => x"00000002",
  2915 => x"00003308",
  2916 => x"000027d3",
  2917 => x"00000002",
  2918 => x"00003326",
  2919 => x"000027d3",
  2920 => x"00000002",
  2921 => x"00003344",
  2922 => x"000027d3",
  2923 => x"00000002",
  2924 => x"00003362",
  2925 => x"000027d3",
  2926 => x"00000002",
  2927 => x"00003380",
  2928 => x"000027d3",
  2929 => x"00000004",
  2930 => x"00002bd8",
  2931 => x"00000000",
  2932 => x"00000000",
  2933 => x"00000000",
  2934 => x"00002994",
  2935 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

