-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80d9",
     9 => x"bc080b0b",
    10 => x"80d9c008",
    11 => x"0b0b80d9",
    12 => x"c4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"d9c40c0b",
    16 => x"0b80d9c0",
    17 => x"0c0b0b80",
    18 => x"d9bc0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d2d4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80d9bc70",
    57 => x"80e4fc27",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a5e3",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80d9",
    65 => x"cc0c9f0b",
    66 => x"80d9d00c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"d9d008ff",
    70 => x"0580d9d0",
    71 => x"0c80d9d0",
    72 => x"088025e8",
    73 => x"3880d9cc",
    74 => x"08ff0580",
    75 => x"d9cc0c80",
    76 => x"d9cc0880",
    77 => x"25d03880",
    78 => x"0b80d9d0",
    79 => x"0c800b80",
    80 => x"d9cc0c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80d9cc08",
   100 => x"25913882",
   101 => x"c82d80d9",
   102 => x"cc08ff05",
   103 => x"80d9cc0c",
   104 => x"838a0480",
   105 => x"d9cc0880",
   106 => x"d9d00853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80d9cc08",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"d9d00881",
   116 => x"0580d9d0",
   117 => x"0c80d9d0",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80d9d0",
   121 => x"0c80d9cc",
   122 => x"08810580",
   123 => x"d9cc0c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480d9",
   128 => x"d0088105",
   129 => x"80d9d00c",
   130 => x"80d9d008",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80d9d0",
   134 => x"0c80d9cc",
   135 => x"08810580",
   136 => x"d9cc0c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"d9d40cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"d9d40c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280d9",
   177 => x"d4088407",
   178 => x"80d9d40c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80d5",
   183 => x"e00c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80d9d4",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80d9",
   208 => x"bc0c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02f8050d",
  1093 => x"028f0580",
  1094 => x"f52d80d5",
  1095 => x"e8085252",
  1096 => x"7080dae9",
  1097 => x"279a3871",
  1098 => x"7181b72d",
  1099 => x"80d5e808",
  1100 => x"810580d5",
  1101 => x"e80c80d5",
  1102 => x"e8085180",
  1103 => x"7181b72d",
  1104 => x"0288050d",
  1105 => x"0402f405",
  1106 => x"0d747084",
  1107 => x"2a708f06",
  1108 => x"80d5e408",
  1109 => x"057080f5",
  1110 => x"2d545153",
  1111 => x"53a2902d",
  1112 => x"728f0680",
  1113 => x"d5e40805",
  1114 => x"7080f52d",
  1115 => x"5253a290",
  1116 => x"2d028c05",
  1117 => x"0d0402f4",
  1118 => x"050d7476",
  1119 => x"54527270",
  1120 => x"81055480",
  1121 => x"f52d5170",
  1122 => x"72708105",
  1123 => x"5481b72d",
  1124 => x"70ec3870",
  1125 => x"7281b72d",
  1126 => x"028c050d",
  1127 => x"0402dc05",
  1128 => x"0d805981",
  1129 => x"0bec0c84",
  1130 => x"0bec0c7a",
  1131 => x"5280d9d8",
  1132 => x"5180c9a2",
  1133 => x"2d80d9bc",
  1134 => x"08792e80",
  1135 => x"f43880d9",
  1136 => x"dc0879ff",
  1137 => x"12565956",
  1138 => x"73792e8b",
  1139 => x"38811874",
  1140 => x"812a5558",
  1141 => x"73f738f7",
  1142 => x"18588159",
  1143 => x"80762580",
  1144 => x"d0387752",
  1145 => x"735184a8",
  1146 => x"2d80dbb4",
  1147 => x"5280d9d8",
  1148 => x"5180cbf6",
  1149 => x"2d80d9bc",
  1150 => x"08802e9b",
  1151 => x"3880dbb4",
  1152 => x"5783fc55",
  1153 => x"76708405",
  1154 => x"5808e80c",
  1155 => x"fc155574",
  1156 => x"8025f138",
  1157 => x"a49f0480",
  1158 => x"d9bc0859",
  1159 => x"84805680",
  1160 => x"d9d85180",
  1161 => x"cbc52dfc",
  1162 => x"80168115",
  1163 => x"5556a3dc",
  1164 => x"0480d9dc",
  1165 => x"08f80c80",
  1166 => x"5186da2d",
  1167 => x"78802e88",
  1168 => x"3880d5ec",
  1169 => x"51a4cc04",
  1170 => x"80d78851",
  1171 => x"add52d78",
  1172 => x"80d9bc0c",
  1173 => x"02a4050d",
  1174 => x"0402f005",
  1175 => x"0d80daa8",
  1176 => x"0b80d5e8",
  1177 => x"0c800b80",
  1178 => x"daa80b81",
  1179 => x"b72d80d7",
  1180 => x"ac0851a2",
  1181 => x"c52dba51",
  1182 => x"a2902d80",
  1183 => x"5480d7ac",
  1184 => x"0814822b",
  1185 => x"f4801108",
  1186 => x"70535153",
  1187 => x"a2c52da0",
  1188 => x"51a2902d",
  1189 => x"72882a51",
  1190 => x"a2c52da0",
  1191 => x"51a2902d",
  1192 => x"72902a51",
  1193 => x"a2c52da0",
  1194 => x"51a2902d",
  1195 => x"72982a51",
  1196 => x"a2c52d81",
  1197 => x"14548174",
  1198 => x"25c33880",
  1199 => x"daa85280",
  1200 => x"d9e451a2",
  1201 => x"f62d80d5",
  1202 => x"ec51add5",
  1203 => x"2d80d7ac",
  1204 => x"08810580",
  1205 => x"d7ac0c02",
  1206 => x"90050d04",
  1207 => x"800b80d7",
  1208 => x"ac0c0402",
  1209 => x"ec050d84",
  1210 => x"0bec0cab",
  1211 => x"922da7c7",
  1212 => x"2d81f92d",
  1213 => x"8353aaf5",
  1214 => x"2d815185",
  1215 => x"8d2dff13",
  1216 => x"53728025",
  1217 => x"f138840b",
  1218 => x"ec0c80d4",
  1219 => x"845186a0",
  1220 => x"2dbfcd2d",
  1221 => x"80d9bc08",
  1222 => x"802e8194",
  1223 => x"38a39d51",
  1224 => x"80d2cb2d",
  1225 => x"80d49c52",
  1226 => x"80d9e451",
  1227 => x"a2f62d80",
  1228 => x"d5ec51ad",
  1229 => x"d52dabb4",
  1230 => x"2da7d32d",
  1231 => x"ade82d80",
  1232 => x"d6800b80",
  1233 => x"f52d80d7",
  1234 => x"f8087081",
  1235 => x"06555654",
  1236 => x"72802e85",
  1237 => x"38738407",
  1238 => x"5474812a",
  1239 => x"70810651",
  1240 => x"5372802e",
  1241 => x"85387382",
  1242 => x"07547482",
  1243 => x"2a708106",
  1244 => x"51537280",
  1245 => x"2e853873",
  1246 => x"81075474",
  1247 => x"832a7081",
  1248 => x"06515372",
  1249 => x"802e8538",
  1250 => x"73880754",
  1251 => x"74842a70",
  1252 => x"81065153",
  1253 => x"72802e85",
  1254 => x"38739007",
  1255 => x"5473fc0c",
  1256 => x"865380d9",
  1257 => x"bc088338",
  1258 => x"845372ec",
  1259 => x"0ca6b904",
  1260 => x"800b80d9",
  1261 => x"bc0c0294",
  1262 => x"050d0471",
  1263 => x"980c04ff",
  1264 => x"b00880d9",
  1265 => x"bc0c0481",
  1266 => x"0bffb00c",
  1267 => x"04800bff",
  1268 => x"b00c0402",
  1269 => x"f4050da8",
  1270 => x"e10480d9",
  1271 => x"bc0881f0",
  1272 => x"2e098106",
  1273 => x"8a38810b",
  1274 => x"80d7f00c",
  1275 => x"a8e10480",
  1276 => x"d9bc0881",
  1277 => x"e02e0981",
  1278 => x"068a3881",
  1279 => x"0b80d7f4",
  1280 => x"0ca8e104",
  1281 => x"80d9bc08",
  1282 => x"5280d7f4",
  1283 => x"08802e89",
  1284 => x"3880d9bc",
  1285 => x"08818005",
  1286 => x"5271842c",
  1287 => x"728f0653",
  1288 => x"5380d7f0",
  1289 => x"08802e9a",
  1290 => x"38728429",
  1291 => x"80d7b005",
  1292 => x"72138171",
  1293 => x"2b700973",
  1294 => x"0806730c",
  1295 => x"515353a8",
  1296 => x"d5047284",
  1297 => x"2980d7b0",
  1298 => x"05721383",
  1299 => x"712b7208",
  1300 => x"07720c53",
  1301 => x"53800b80",
  1302 => x"d7f40c80",
  1303 => x"0b80d7f0",
  1304 => x"0c80daec",
  1305 => x"51a9e82d",
  1306 => x"80d9bc08",
  1307 => x"ff24feea",
  1308 => x"38800b80",
  1309 => x"d9bc0c02",
  1310 => x"8c050d04",
  1311 => x"02f8050d",
  1312 => x"80d7b052",
  1313 => x"8f518072",
  1314 => x"70840554",
  1315 => x"0cff1151",
  1316 => x"708025f2",
  1317 => x"38028805",
  1318 => x"0d0402f0",
  1319 => x"050d7551",
  1320 => x"a7cd2d70",
  1321 => x"822cfc06",
  1322 => x"80d7b011",
  1323 => x"72109e06",
  1324 => x"71087072",
  1325 => x"2a708306",
  1326 => x"82742b70",
  1327 => x"09740676",
  1328 => x"0c545156",
  1329 => x"57535153",
  1330 => x"a7c72d71",
  1331 => x"80d9bc0c",
  1332 => x"0290050d",
  1333 => x"0402fc05",
  1334 => x"0d725180",
  1335 => x"710c800b",
  1336 => x"84120c02",
  1337 => x"84050d04",
  1338 => x"02f0050d",
  1339 => x"75700884",
  1340 => x"12085353",
  1341 => x"53ff5471",
  1342 => x"712ea838",
  1343 => x"a7cd2d84",
  1344 => x"13087084",
  1345 => x"29148811",
  1346 => x"70087081",
  1347 => x"ff068418",
  1348 => x"08811187",
  1349 => x"06841a0c",
  1350 => x"53515551",
  1351 => x"5151a7c7",
  1352 => x"2d715473",
  1353 => x"80d9bc0c",
  1354 => x"0290050d",
  1355 => x"0402f805",
  1356 => x"0da7cd2d",
  1357 => x"e008708b",
  1358 => x"2a708106",
  1359 => x"51525270",
  1360 => x"802ea138",
  1361 => x"80daec08",
  1362 => x"70842980",
  1363 => x"daf40573",
  1364 => x"81ff0671",
  1365 => x"0c515180",
  1366 => x"daec0881",
  1367 => x"11870680",
  1368 => x"daec0c51",
  1369 => x"800b80db",
  1370 => x"940ca7bf",
  1371 => x"2da7c72d",
  1372 => x"0288050d",
  1373 => x"0402fc05",
  1374 => x"0da7cd2d",
  1375 => x"810b80db",
  1376 => x"940ca7c7",
  1377 => x"2d80db94",
  1378 => x"085170f9",
  1379 => x"38028405",
  1380 => x"0d0402fc",
  1381 => x"050d80da",
  1382 => x"ec51a9d5",
  1383 => x"2da8fc2d",
  1384 => x"aaad51a7",
  1385 => x"bb2d0284",
  1386 => x"050d0480",
  1387 => x"dba00880",
  1388 => x"d9bc0c04",
  1389 => x"02fc050d",
  1390 => x"810b80d7",
  1391 => x"fc0c8151",
  1392 => x"858d2d02",
  1393 => x"84050d04",
  1394 => x"02fc050d",
  1395 => x"abd204a7",
  1396 => x"d32d80f6",
  1397 => x"51a99a2d",
  1398 => x"80d9bc08",
  1399 => x"f23880da",
  1400 => x"51a99a2d",
  1401 => x"80d9bc08",
  1402 => x"e63880d9",
  1403 => x"bc0880d7",
  1404 => x"fc0c80d9",
  1405 => x"bc085185",
  1406 => x"8d2d0284",
  1407 => x"050d0402",
  1408 => x"ec050d76",
  1409 => x"54805287",
  1410 => x"0b881580",
  1411 => x"f52d5653",
  1412 => x"74722483",
  1413 => x"38a05372",
  1414 => x"5183842d",
  1415 => x"81128b15",
  1416 => x"80f52d54",
  1417 => x"52727225",
  1418 => x"de380294",
  1419 => x"050d0402",
  1420 => x"f0050d80",
  1421 => x"dba00854",
  1422 => x"81f92d80",
  1423 => x"0b80dba4",
  1424 => x"0c730880",
  1425 => x"2e818938",
  1426 => x"820b80d9",
  1427 => x"d00c80db",
  1428 => x"a4088f06",
  1429 => x"80d9cc0c",
  1430 => x"73085271",
  1431 => x"832e9638",
  1432 => x"71832689",
  1433 => x"3871812e",
  1434 => x"b038adb9",
  1435 => x"0471852e",
  1436 => x"a038adb9",
  1437 => x"04881480",
  1438 => x"f52d8415",
  1439 => x"0880d4ac",
  1440 => x"53545286",
  1441 => x"a02d7184",
  1442 => x"29137008",
  1443 => x"5252adbd",
  1444 => x"047351ab",
  1445 => x"ff2dadb9",
  1446 => x"0480d7f8",
  1447 => x"08881508",
  1448 => x"2c708106",
  1449 => x"51527180",
  1450 => x"2e883880",
  1451 => x"d4b051ad",
  1452 => x"b60480d4",
  1453 => x"b45186a0",
  1454 => x"2d841408",
  1455 => x"5186a02d",
  1456 => x"80dba408",
  1457 => x"810580db",
  1458 => x"a40c8c14",
  1459 => x"54acc104",
  1460 => x"0290050d",
  1461 => x"047180db",
  1462 => x"a00cacaf",
  1463 => x"2d80dba4",
  1464 => x"08ff0580",
  1465 => x"dba80c04",
  1466 => x"02e8050d",
  1467 => x"80dba008",
  1468 => x"80dbac08",
  1469 => x"575580f6",
  1470 => x"51a99a2d",
  1471 => x"80d9bc08",
  1472 => x"812a7081",
  1473 => x"06515271",
  1474 => x"802ea438",
  1475 => x"ae9204a7",
  1476 => x"d32d80f6",
  1477 => x"51a99a2d",
  1478 => x"80d9bc08",
  1479 => x"f23880d7",
  1480 => x"fc088132",
  1481 => x"7080d7fc",
  1482 => x"0c705252",
  1483 => x"858d2d80",
  1484 => x"0b80db98",
  1485 => x"0c800b80",
  1486 => x"db9c0c80",
  1487 => x"d7fc0883",
  1488 => x"8d3880da",
  1489 => x"51a99a2d",
  1490 => x"80d9bc08",
  1491 => x"802e8c38",
  1492 => x"80db9808",
  1493 => x"81800780",
  1494 => x"db980c80",
  1495 => x"d951a99a",
  1496 => x"2d80d9bc",
  1497 => x"08802e8c",
  1498 => x"3880db98",
  1499 => x"0880c007",
  1500 => x"80db980c",
  1501 => x"819451a9",
  1502 => x"9a2d80d9",
  1503 => x"bc08802e",
  1504 => x"8b3880db",
  1505 => x"98089007",
  1506 => x"80db980c",
  1507 => x"819151a9",
  1508 => x"9a2d80d9",
  1509 => x"bc08802e",
  1510 => x"8b3880db",
  1511 => x"9808a007",
  1512 => x"80db980c",
  1513 => x"81f551a9",
  1514 => x"9a2d80d9",
  1515 => x"bc08802e",
  1516 => x"8b3880db",
  1517 => x"98088107",
  1518 => x"80db980c",
  1519 => x"81f251a9",
  1520 => x"9a2d80d9",
  1521 => x"bc08802e",
  1522 => x"8b3880db",
  1523 => x"98088207",
  1524 => x"80db980c",
  1525 => x"81eb51a9",
  1526 => x"9a2d80d9",
  1527 => x"bc08802e",
  1528 => x"8b3880db",
  1529 => x"98088407",
  1530 => x"80db980c",
  1531 => x"81f451a9",
  1532 => x"9a2d80d9",
  1533 => x"bc08802e",
  1534 => x"8b3880db",
  1535 => x"98088807",
  1536 => x"80db980c",
  1537 => x"80d851a9",
  1538 => x"9a2d80d9",
  1539 => x"bc08802e",
  1540 => x"8c3880db",
  1541 => x"9c088180",
  1542 => x"0780db9c",
  1543 => x"0c9251a9",
  1544 => x"9a2d80d9",
  1545 => x"bc08802e",
  1546 => x"8c3880db",
  1547 => x"9c0880c0",
  1548 => x"0780db9c",
  1549 => x"0c9451a9",
  1550 => x"9a2d80d9",
  1551 => x"bc08802e",
  1552 => x"8b3880db",
  1553 => x"9c089007",
  1554 => x"80db9c0c",
  1555 => x"9151a99a",
  1556 => x"2d80d9bc",
  1557 => x"08802e8b",
  1558 => x"3880db9c",
  1559 => x"08a00780",
  1560 => x"db9c0c9d",
  1561 => x"51a99a2d",
  1562 => x"80d9bc08",
  1563 => x"802e8b38",
  1564 => x"80db9c08",
  1565 => x"810780db",
  1566 => x"9c0c9b51",
  1567 => x"a99a2d80",
  1568 => x"d9bc0880",
  1569 => x"2e8b3880",
  1570 => x"db9c0882",
  1571 => x"0780db9c",
  1572 => x"0c9c51a9",
  1573 => x"9a2d80d9",
  1574 => x"bc08802e",
  1575 => x"8b3880db",
  1576 => x"9c088407",
  1577 => x"80db9c0c",
  1578 => x"a351a99a",
  1579 => x"2d80d9bc",
  1580 => x"08802e8b",
  1581 => x"3880db9c",
  1582 => x"08880780",
  1583 => x"db9c0c81",
  1584 => x"fd51a99a",
  1585 => x"2d81fa51",
  1586 => x"a99a2db7",
  1587 => x"a30481f5",
  1588 => x"51a99a2d",
  1589 => x"80d9bc08",
  1590 => x"812a7081",
  1591 => x"06515271",
  1592 => x"802eb338",
  1593 => x"80dba808",
  1594 => x"5271802e",
  1595 => x"8a38ff12",
  1596 => x"80dba80c",
  1597 => x"b2960480",
  1598 => x"dba40810",
  1599 => x"80dba408",
  1600 => x"05708429",
  1601 => x"16515288",
  1602 => x"1208802e",
  1603 => x"8938ff51",
  1604 => x"88120852",
  1605 => x"712d81f2",
  1606 => x"51a99a2d",
  1607 => x"80d9bc08",
  1608 => x"812a7081",
  1609 => x"06515271",
  1610 => x"802eb438",
  1611 => x"80dba408",
  1612 => x"ff1180db",
  1613 => x"a8085653",
  1614 => x"53737225",
  1615 => x"8a388114",
  1616 => x"80dba80c",
  1617 => x"b2df0472",
  1618 => x"10137084",
  1619 => x"29165152",
  1620 => x"88120880",
  1621 => x"2e8938fe",
  1622 => x"51881208",
  1623 => x"52712d81",
  1624 => x"fd51a99a",
  1625 => x"2d80d9bc",
  1626 => x"08812a70",
  1627 => x"81065152",
  1628 => x"71802eb1",
  1629 => x"3880dba8",
  1630 => x"08802e8a",
  1631 => x"38800b80",
  1632 => x"dba80cb3",
  1633 => x"a50480db",
  1634 => x"a4081080",
  1635 => x"dba40805",
  1636 => x"70842916",
  1637 => x"51528812",
  1638 => x"08802e89",
  1639 => x"38fd5188",
  1640 => x"12085271",
  1641 => x"2d81fa51",
  1642 => x"a99a2d80",
  1643 => x"d9bc0881",
  1644 => x"2a708106",
  1645 => x"51527180",
  1646 => x"2eb13880",
  1647 => x"dba408ff",
  1648 => x"11545280",
  1649 => x"dba80873",
  1650 => x"25893872",
  1651 => x"80dba80c",
  1652 => x"b3eb0471",
  1653 => x"10127084",
  1654 => x"29165152",
  1655 => x"88120880",
  1656 => x"2e8938fc",
  1657 => x"51881208",
  1658 => x"52712d80",
  1659 => x"dba80870",
  1660 => x"53547380",
  1661 => x"2e8a388c",
  1662 => x"15ff1555",
  1663 => x"55b3f204",
  1664 => x"820b80d9",
  1665 => x"d00c718f",
  1666 => x"0680d9cc",
  1667 => x"0c81eb51",
  1668 => x"a99a2d80",
  1669 => x"d9bc0881",
  1670 => x"2a708106",
  1671 => x"51527180",
  1672 => x"2ead3874",
  1673 => x"08852e09",
  1674 => x"8106a438",
  1675 => x"881580f5",
  1676 => x"2dff0552",
  1677 => x"71881681",
  1678 => x"b72d7198",
  1679 => x"2b527180",
  1680 => x"25883880",
  1681 => x"0b881681",
  1682 => x"b72d7451",
  1683 => x"abff2d81",
  1684 => x"f451a99a",
  1685 => x"2d80d9bc",
  1686 => x"08812a70",
  1687 => x"81065152",
  1688 => x"71802eb3",
  1689 => x"38740885",
  1690 => x"2e098106",
  1691 => x"aa388815",
  1692 => x"80f52d81",
  1693 => x"05527188",
  1694 => x"1681b72d",
  1695 => x"7181ff06",
  1696 => x"8b1680f5",
  1697 => x"2d545272",
  1698 => x"72278738",
  1699 => x"72881681",
  1700 => x"b72d7451",
  1701 => x"abff2d80",
  1702 => x"da51a99a",
  1703 => x"2d80d9bc",
  1704 => x"08812a70",
  1705 => x"81065152",
  1706 => x"71802e81",
  1707 => x"ad3880db",
  1708 => x"a00880db",
  1709 => x"a8085553",
  1710 => x"73802e8a",
  1711 => x"388c13ff",
  1712 => x"155553b5",
  1713 => x"b8047208",
  1714 => x"5271822e",
  1715 => x"a6387182",
  1716 => x"26893871",
  1717 => x"812eaa38",
  1718 => x"b6da0471",
  1719 => x"832eb438",
  1720 => x"71842e09",
  1721 => x"810680f2",
  1722 => x"38881308",
  1723 => x"51add52d",
  1724 => x"b6da0480",
  1725 => x"dba80851",
  1726 => x"88130852",
  1727 => x"712db6da",
  1728 => x"04810b88",
  1729 => x"14082b80",
  1730 => x"d7f80832",
  1731 => x"80d7f80c",
  1732 => x"b6ae0488",
  1733 => x"1380f52d",
  1734 => x"81058b14",
  1735 => x"80f52d53",
  1736 => x"54717424",
  1737 => x"83388054",
  1738 => x"73881481",
  1739 => x"b72dacaf",
  1740 => x"2db6da04",
  1741 => x"7508802e",
  1742 => x"a4387508",
  1743 => x"51a99a2d",
  1744 => x"80d9bc08",
  1745 => x"81065271",
  1746 => x"802e8c38",
  1747 => x"80dba808",
  1748 => x"51841608",
  1749 => x"52712d88",
  1750 => x"165675d8",
  1751 => x"38805480",
  1752 => x"0b80d9d0",
  1753 => x"0c738f06",
  1754 => x"80d9cc0c",
  1755 => x"a0527380",
  1756 => x"dba8082e",
  1757 => x"09810699",
  1758 => x"3880dba4",
  1759 => x"08ff0574",
  1760 => x"32700981",
  1761 => x"05707207",
  1762 => x"9f2a9171",
  1763 => x"31515153",
  1764 => x"53715183",
  1765 => x"842d8114",
  1766 => x"548e7425",
  1767 => x"c23880d7",
  1768 => x"fc085271",
  1769 => x"80d9bc0c",
  1770 => x"0298050d",
  1771 => x"0402f405",
  1772 => x"0dd45281",
  1773 => x"ff720c71",
  1774 => x"085381ff",
  1775 => x"720c7288",
  1776 => x"2b83fe80",
  1777 => x"06720870",
  1778 => x"81ff0651",
  1779 => x"525381ff",
  1780 => x"720c7271",
  1781 => x"07882b72",
  1782 => x"087081ff",
  1783 => x"06515253",
  1784 => x"81ff720c",
  1785 => x"72710788",
  1786 => x"2b720870",
  1787 => x"81ff0672",
  1788 => x"0780d9bc",
  1789 => x"0c525302",
  1790 => x"8c050d04",
  1791 => x"02f4050d",
  1792 => x"74767181",
  1793 => x"ff06d40c",
  1794 => x"535380db",
  1795 => x"b0088538",
  1796 => x"71892b52",
  1797 => x"71982ad4",
  1798 => x"0c71902a",
  1799 => x"7081ff06",
  1800 => x"d40c5171",
  1801 => x"882a7081",
  1802 => x"ff06d40c",
  1803 => x"517181ff",
  1804 => x"06d40c72",
  1805 => x"902a7081",
  1806 => x"ff06d40c",
  1807 => x"51d40870",
  1808 => x"81ff0651",
  1809 => x"5182b8bf",
  1810 => x"527081ff",
  1811 => x"2e098106",
  1812 => x"943881ff",
  1813 => x"0bd40cd4",
  1814 => x"087081ff",
  1815 => x"06ff1454",
  1816 => x"515171e5",
  1817 => x"387080d9",
  1818 => x"bc0c028c",
  1819 => x"050d0402",
  1820 => x"fc050d81",
  1821 => x"c75181ff",
  1822 => x"0bd40cff",
  1823 => x"11517080",
  1824 => x"25f43802",
  1825 => x"84050d04",
  1826 => x"02f4050d",
  1827 => x"81ff0bd4",
  1828 => x"0c935380",
  1829 => x"5287fc80",
  1830 => x"c151b7fc",
  1831 => x"2d80d9bc",
  1832 => x"088b3881",
  1833 => x"ff0bd40c",
  1834 => x"8153b9b6",
  1835 => x"04b8ef2d",
  1836 => x"ff135372",
  1837 => x"de387280",
  1838 => x"d9bc0c02",
  1839 => x"8c050d04",
  1840 => x"02ec050d",
  1841 => x"810b80db",
  1842 => x"b00c8454",
  1843 => x"d008708f",
  1844 => x"2a708106",
  1845 => x"51515372",
  1846 => x"f33872d0",
  1847 => x"0cb8ef2d",
  1848 => x"80d4b851",
  1849 => x"86a02dd0",
  1850 => x"08708f2a",
  1851 => x"70810651",
  1852 => x"515372f3",
  1853 => x"38810bd0",
  1854 => x"0cb15380",
  1855 => x"5284d480",
  1856 => x"c051b7fc",
  1857 => x"2d80d9bc",
  1858 => x"08812e93",
  1859 => x"3872822e",
  1860 => x"bf38ff13",
  1861 => x"5372e438",
  1862 => x"ff145473",
  1863 => x"ffae38b8",
  1864 => x"ef2d83aa",
  1865 => x"52849c80",
  1866 => x"c851b7fc",
  1867 => x"2d80d9bc",
  1868 => x"08812e09",
  1869 => x"81069338",
  1870 => x"b7ad2d80",
  1871 => x"d9bc0883",
  1872 => x"ffff0653",
  1873 => x"7283aa2e",
  1874 => x"9f38b988",
  1875 => x"2dbae304",
  1876 => x"80d4c451",
  1877 => x"86a02d80",
  1878 => x"53bcb804",
  1879 => x"80d4dc51",
  1880 => x"86a02d80",
  1881 => x"54bc8904",
  1882 => x"81ff0bd4",
  1883 => x"0cb154b8",
  1884 => x"ef2d8fcf",
  1885 => x"53805287",
  1886 => x"fc80f751",
  1887 => x"b7fc2d80",
  1888 => x"d9bc0855",
  1889 => x"80d9bc08",
  1890 => x"812e0981",
  1891 => x"069c3881",
  1892 => x"ff0bd40c",
  1893 => x"820a5284",
  1894 => x"9c80e951",
  1895 => x"b7fc2d80",
  1896 => x"d9bc0880",
  1897 => x"2e8d38b8",
  1898 => x"ef2dff13",
  1899 => x"5372c638",
  1900 => x"bbfc0481",
  1901 => x"ff0bd40c",
  1902 => x"80d9bc08",
  1903 => x"5287fc80",
  1904 => x"fa51b7fc",
  1905 => x"2d80d9bc",
  1906 => x"08b23881",
  1907 => x"ff0bd40c",
  1908 => x"d4085381",
  1909 => x"ff0bd40c",
  1910 => x"81ff0bd4",
  1911 => x"0c81ff0b",
  1912 => x"d40c81ff",
  1913 => x"0bd40c72",
  1914 => x"862a7081",
  1915 => x"06765651",
  1916 => x"53729638",
  1917 => x"80d9bc08",
  1918 => x"54bc8904",
  1919 => x"73822efe",
  1920 => x"db38ff14",
  1921 => x"5473fee7",
  1922 => x"387380db",
  1923 => x"b00c738b",
  1924 => x"38815287",
  1925 => x"fc80d051",
  1926 => x"b7fc2d81",
  1927 => x"ff0bd40c",
  1928 => x"d008708f",
  1929 => x"2a708106",
  1930 => x"51515372",
  1931 => x"f33872d0",
  1932 => x"0c81ff0b",
  1933 => x"d40c8153",
  1934 => x"7280d9bc",
  1935 => x"0c029405",
  1936 => x"0d0402e8",
  1937 => x"050d7855",
  1938 => x"805681ff",
  1939 => x"0bd40cd0",
  1940 => x"08708f2a",
  1941 => x"70810651",
  1942 => x"515372f3",
  1943 => x"3882810b",
  1944 => x"d00c81ff",
  1945 => x"0bd40c77",
  1946 => x"5287fc80",
  1947 => x"d151b7fc",
  1948 => x"2d80dbc6",
  1949 => x"df5480d9",
  1950 => x"bc08802e",
  1951 => x"8b3880d4",
  1952 => x"fc5186a0",
  1953 => x"2dbddc04",
  1954 => x"81ff0bd4",
  1955 => x"0cd40870",
  1956 => x"81ff0651",
  1957 => x"537281fe",
  1958 => x"2e098106",
  1959 => x"9e3880ff",
  1960 => x"53b7ad2d",
  1961 => x"80d9bc08",
  1962 => x"75708405",
  1963 => x"570cff13",
  1964 => x"53728025",
  1965 => x"ec388156",
  1966 => x"bdc104ff",
  1967 => x"145473c8",
  1968 => x"3881ff0b",
  1969 => x"d40c81ff",
  1970 => x"0bd40cd0",
  1971 => x"08708f2a",
  1972 => x"70810651",
  1973 => x"515372f3",
  1974 => x"3872d00c",
  1975 => x"7580d9bc",
  1976 => x"0c029805",
  1977 => x"0d0402e8",
  1978 => x"050d7779",
  1979 => x"7b585555",
  1980 => x"80537276",
  1981 => x"25a33874",
  1982 => x"70810556",
  1983 => x"80f52d74",
  1984 => x"70810556",
  1985 => x"80f52d52",
  1986 => x"5271712e",
  1987 => x"86388151",
  1988 => x"be9b0481",
  1989 => x"1353bdf2",
  1990 => x"04805170",
  1991 => x"80d9bc0c",
  1992 => x"0298050d",
  1993 => x"0402ec05",
  1994 => x"0d765574",
  1995 => x"802e80c4",
  1996 => x"389a1580",
  1997 => x"e02d5180",
  1998 => x"ccd02d80",
  1999 => x"d9bc0880",
  2000 => x"d9bc0880",
  2001 => x"e1e40c80",
  2002 => x"d9bc0854",
  2003 => x"5480e1c0",
  2004 => x"08802e9b",
  2005 => x"38941580",
  2006 => x"e02d5180",
  2007 => x"ccd02d80",
  2008 => x"d9bc0890",
  2009 => x"2b83fff0",
  2010 => x"0a067075",
  2011 => x"07515372",
  2012 => x"80e1e40c",
  2013 => x"80e1e408",
  2014 => x"5372802e",
  2015 => x"9d3880e1",
  2016 => x"b808fe14",
  2017 => x"712980e1",
  2018 => x"cc080580",
  2019 => x"e1e80c70",
  2020 => x"842b80e1",
  2021 => x"c40c54bf",
  2022 => x"c80480e1",
  2023 => x"d00880e1",
  2024 => x"e40c80e1",
  2025 => x"d40880e1",
  2026 => x"e80c80e1",
  2027 => x"c008802e",
  2028 => x"8b3880e1",
  2029 => x"b808842b",
  2030 => x"53bfc304",
  2031 => x"80e1d808",
  2032 => x"842b5372",
  2033 => x"80e1c40c",
  2034 => x"0294050d",
  2035 => x"0402d805",
  2036 => x"0d800b80",
  2037 => x"e1c00c84",
  2038 => x"54b9c02d",
  2039 => x"80d9bc08",
  2040 => x"802e9838",
  2041 => x"80dbb452",
  2042 => x"8051bcc2",
  2043 => x"2d80d9bc",
  2044 => x"08802e87",
  2045 => x"38fe5480",
  2046 => x"c08304ff",
  2047 => x"14547380",
  2048 => x"24d73873",
  2049 => x"8e3880d5",
  2050 => x"8c5186a0",
  2051 => x"2d735580",
  2052 => x"c5e00480",
  2053 => x"56810b80",
  2054 => x"e1ec0c88",
  2055 => x"5380d5a0",
  2056 => x"5280dbea",
  2057 => x"51bde62d",
  2058 => x"80d9bc08",
  2059 => x"762e0981",
  2060 => x"06893880",
  2061 => x"d9bc0880",
  2062 => x"e1ec0c88",
  2063 => x"5380d5ac",
  2064 => x"5280dc86",
  2065 => x"51bde62d",
  2066 => x"80d9bc08",
  2067 => x"893880d9",
  2068 => x"bc0880e1",
  2069 => x"ec0c80e1",
  2070 => x"ec08802e",
  2071 => x"81843880",
  2072 => x"defa0b80",
  2073 => x"f52d80de",
  2074 => x"fb0b80f5",
  2075 => x"2d71982b",
  2076 => x"71902b07",
  2077 => x"80defc0b",
  2078 => x"80f52d70",
  2079 => x"882b7207",
  2080 => x"80defd0b",
  2081 => x"80f52d71",
  2082 => x"0780dfb2",
  2083 => x"0b80f52d",
  2084 => x"80dfb30b",
  2085 => x"80f52d71",
  2086 => x"882b0753",
  2087 => x"5f54525a",
  2088 => x"56575573",
  2089 => x"81abaa2e",
  2090 => x"09810690",
  2091 => x"38755180",
  2092 => x"cc9f2d80",
  2093 => x"d9bc0856",
  2094 => x"80c1cb04",
  2095 => x"7382d4d5",
  2096 => x"2e893880",
  2097 => x"d5b85180",
  2098 => x"c2980480",
  2099 => x"dbb45275",
  2100 => x"51bcc22d",
  2101 => x"80d9bc08",
  2102 => x"5580d9bc",
  2103 => x"08802e83",
  2104 => x"ff388853",
  2105 => x"80d5ac52",
  2106 => x"80dc8651",
  2107 => x"bde62d80",
  2108 => x"d9bc088b",
  2109 => x"38810b80",
  2110 => x"e1c00c80",
  2111 => x"c29f0488",
  2112 => x"5380d5a0",
  2113 => x"5280dbea",
  2114 => x"51bde62d",
  2115 => x"80d9bc08",
  2116 => x"802e8c38",
  2117 => x"80d5cc51",
  2118 => x"86a02d80",
  2119 => x"c2fe0480",
  2120 => x"dfb20b80",
  2121 => x"f52d5473",
  2122 => x"80d52e09",
  2123 => x"810680ce",
  2124 => x"3880dfb3",
  2125 => x"0b80f52d",
  2126 => x"547381aa",
  2127 => x"2e098106",
  2128 => x"bd38800b",
  2129 => x"80dbb40b",
  2130 => x"80f52d56",
  2131 => x"547481e9",
  2132 => x"2e833881",
  2133 => x"547481eb",
  2134 => x"2e8c3880",
  2135 => x"5573752e",
  2136 => x"09810682",
  2137 => x"fb3880db",
  2138 => x"bf0b80f5",
  2139 => x"2d55748e",
  2140 => x"3880dbc0",
  2141 => x"0b80f52d",
  2142 => x"5473822e",
  2143 => x"87388055",
  2144 => x"80c5e004",
  2145 => x"80dbc10b",
  2146 => x"80f52d70",
  2147 => x"80e1b80c",
  2148 => x"ff0580e1",
  2149 => x"bc0c80db",
  2150 => x"c20b80f5",
  2151 => x"2d80dbc3",
  2152 => x"0b80f52d",
  2153 => x"58760577",
  2154 => x"82802905",
  2155 => x"7080e1c8",
  2156 => x"0c80dbc4",
  2157 => x"0b80f52d",
  2158 => x"7080e1dc",
  2159 => x"0c80e1c0",
  2160 => x"08595758",
  2161 => x"76802e81",
  2162 => x"b8388853",
  2163 => x"80d5ac52",
  2164 => x"80dc8651",
  2165 => x"bde62d80",
  2166 => x"d9bc0882",
  2167 => x"833880e1",
  2168 => x"b8087084",
  2169 => x"2b80e1c4",
  2170 => x"0c7080e1",
  2171 => x"d80c80db",
  2172 => x"d90b80f5",
  2173 => x"2d80dbd8",
  2174 => x"0b80f52d",
  2175 => x"71828029",
  2176 => x"0580dbda",
  2177 => x"0b80f52d",
  2178 => x"70848080",
  2179 => x"291280db",
  2180 => x"db0b80f5",
  2181 => x"2d708180",
  2182 => x"0a291270",
  2183 => x"80e1e00c",
  2184 => x"80e1dc08",
  2185 => x"712980e1",
  2186 => x"c8080570",
  2187 => x"80e1cc0c",
  2188 => x"80dbe10b",
  2189 => x"80f52d80",
  2190 => x"dbe00b80",
  2191 => x"f52d7182",
  2192 => x"80290580",
  2193 => x"dbe20b80",
  2194 => x"f52d7084",
  2195 => x"80802912",
  2196 => x"80dbe30b",
  2197 => x"80f52d70",
  2198 => x"982b81f0",
  2199 => x"0a067205",
  2200 => x"7080e1d0",
  2201 => x"0cfe117e",
  2202 => x"29770580",
  2203 => x"e1d40c52",
  2204 => x"59524354",
  2205 => x"5e515259",
  2206 => x"525d5759",
  2207 => x"5780c5d9",
  2208 => x"0480dbc6",
  2209 => x"0b80f52d",
  2210 => x"80dbc50b",
  2211 => x"80f52d71",
  2212 => x"82802905",
  2213 => x"7080e1c4",
  2214 => x"0c70a029",
  2215 => x"83ff0570",
  2216 => x"892a7080",
  2217 => x"e1d80c80",
  2218 => x"dbcb0b80",
  2219 => x"f52d80db",
  2220 => x"ca0b80f5",
  2221 => x"2d718280",
  2222 => x"29057080",
  2223 => x"e1e00c7b",
  2224 => x"71291e70",
  2225 => x"80e1d40c",
  2226 => x"7d80e1d0",
  2227 => x"0c730580",
  2228 => x"e1cc0c55",
  2229 => x"5e515155",
  2230 => x"558051be",
  2231 => x"a52d8155",
  2232 => x"7480d9bc",
  2233 => x"0c02a805",
  2234 => x"0d0402ec",
  2235 => x"050d7670",
  2236 => x"872c7180",
  2237 => x"ff065556",
  2238 => x"5480e1c0",
  2239 => x"088a3873",
  2240 => x"882c7481",
  2241 => x"ff065455",
  2242 => x"80dbb452",
  2243 => x"80e1c808",
  2244 => x"1551bcc2",
  2245 => x"2d80d9bc",
  2246 => x"085480d9",
  2247 => x"bc08802e",
  2248 => x"bb3880e1",
  2249 => x"c008802e",
  2250 => x"9c387284",
  2251 => x"2980dbb4",
  2252 => x"05700852",
  2253 => x"5380cc9f",
  2254 => x"2d80d9bc",
  2255 => x"08f00a06",
  2256 => x"5380c6da",
  2257 => x"04721080",
  2258 => x"dbb40570",
  2259 => x"80e02d52",
  2260 => x"5380ccd0",
  2261 => x"2d80d9bc",
  2262 => x"08537254",
  2263 => x"7380d9bc",
  2264 => x"0c029405",
  2265 => x"0d0402e0",
  2266 => x"050d7970",
  2267 => x"842c80e1",
  2268 => x"e8080571",
  2269 => x"8f065255",
  2270 => x"53728a38",
  2271 => x"80dbb452",
  2272 => x"7351bcc2",
  2273 => x"2d72a029",
  2274 => x"80dbb405",
  2275 => x"54807480",
  2276 => x"f52d5653",
  2277 => x"74732e83",
  2278 => x"38815374",
  2279 => x"81e52e81",
  2280 => x"f5388170",
  2281 => x"74065458",
  2282 => x"72802e81",
  2283 => x"e9388b14",
  2284 => x"80f52d70",
  2285 => x"832a7906",
  2286 => x"5856769c",
  2287 => x"3880d880",
  2288 => x"08537289",
  2289 => x"387280df",
  2290 => x"b40b81b7",
  2291 => x"2d7680d8",
  2292 => x"800c7353",
  2293 => x"80c99804",
  2294 => x"758f2e09",
  2295 => x"810681b6",
  2296 => x"38749f06",
  2297 => x"8d2980df",
  2298 => x"a7115153",
  2299 => x"811480f5",
  2300 => x"2d737081",
  2301 => x"055581b7",
  2302 => x"2d831480",
  2303 => x"f52d7370",
  2304 => x"81055581",
  2305 => x"b72d8514",
  2306 => x"80f52d73",
  2307 => x"70810555",
  2308 => x"81b72d87",
  2309 => x"1480f52d",
  2310 => x"73708105",
  2311 => x"5581b72d",
  2312 => x"891480f5",
  2313 => x"2d737081",
  2314 => x"055581b7",
  2315 => x"2d8e1480",
  2316 => x"f52d7370",
  2317 => x"81055581",
  2318 => x"b72d9014",
  2319 => x"80f52d73",
  2320 => x"70810555",
  2321 => x"81b72d92",
  2322 => x"1480f52d",
  2323 => x"73708105",
  2324 => x"5581b72d",
  2325 => x"941480f5",
  2326 => x"2d737081",
  2327 => x"055581b7",
  2328 => x"2d961480",
  2329 => x"f52d7370",
  2330 => x"81055581",
  2331 => x"b72d9814",
  2332 => x"80f52d73",
  2333 => x"70810555",
  2334 => x"81b72d9c",
  2335 => x"1480f52d",
  2336 => x"73708105",
  2337 => x"5581b72d",
  2338 => x"9e1480f5",
  2339 => x"2d7381b7",
  2340 => x"2d7780d8",
  2341 => x"800c8053",
  2342 => x"7280d9bc",
  2343 => x"0c02a005",
  2344 => x"0d0402cc",
  2345 => x"050d7e60",
  2346 => x"5e5a800b",
  2347 => x"80e1e408",
  2348 => x"80e1e808",
  2349 => x"595c5680",
  2350 => x"5880e1c4",
  2351 => x"08782e81",
  2352 => x"bc38778f",
  2353 => x"06a01757",
  2354 => x"54739138",
  2355 => x"80dbb452",
  2356 => x"76518117",
  2357 => x"57bcc22d",
  2358 => x"80dbb456",
  2359 => x"807680f5",
  2360 => x"2d565474",
  2361 => x"742e8338",
  2362 => x"81547481",
  2363 => x"e52e8181",
  2364 => x"38817075",
  2365 => x"06555c73",
  2366 => x"802e80f5",
  2367 => x"388b1680",
  2368 => x"f52d9806",
  2369 => x"597880e9",
  2370 => x"388b537c",
  2371 => x"527551bd",
  2372 => x"e62d80d9",
  2373 => x"bc0880d9",
  2374 => x"389c1608",
  2375 => x"5180cc9f",
  2376 => x"2d80d9bc",
  2377 => x"08841b0c",
  2378 => x"9a1680e0",
  2379 => x"2d5180cc",
  2380 => x"d02d80d9",
  2381 => x"bc0880d9",
  2382 => x"bc08881c",
  2383 => x"0c80d9bc",
  2384 => x"08555580",
  2385 => x"e1c00880",
  2386 => x"2e9a3894",
  2387 => x"1680e02d",
  2388 => x"5180ccd0",
  2389 => x"2d80d9bc",
  2390 => x"08902b83",
  2391 => x"fff00a06",
  2392 => x"70165154",
  2393 => x"73881b0c",
  2394 => x"787a0c7b",
  2395 => x"5480cbbb",
  2396 => x"04811858",
  2397 => x"80e1c408",
  2398 => x"7826fec6",
  2399 => x"3880e1c0",
  2400 => x"08802eb5",
  2401 => x"387a5180",
  2402 => x"c5ea2d80",
  2403 => x"d9bc0880",
  2404 => x"d9bc0880",
  2405 => x"fffffff8",
  2406 => x"06555b73",
  2407 => x"80ffffff",
  2408 => x"f82e9638",
  2409 => x"80d9bc08",
  2410 => x"fe0580e1",
  2411 => x"b8082980",
  2412 => x"e1cc0805",
  2413 => x"5780c9b7",
  2414 => x"04805473",
  2415 => x"80d9bc0c",
  2416 => x"02b4050d",
  2417 => x"0402f405",
  2418 => x"0d747008",
  2419 => x"8105710c",
  2420 => x"700880e1",
  2421 => x"bc080653",
  2422 => x"53719038",
  2423 => x"88130851",
  2424 => x"80c5ea2d",
  2425 => x"80d9bc08",
  2426 => x"88140c81",
  2427 => x"0b80d9bc",
  2428 => x"0c028c05",
  2429 => x"0d0402f0",
  2430 => x"050d7588",
  2431 => x"1108fe05",
  2432 => x"80e1b808",
  2433 => x"2980e1cc",
  2434 => x"08117208",
  2435 => x"80e1bc08",
  2436 => x"06057955",
  2437 => x"535454bc",
  2438 => x"c22d0290",
  2439 => x"050d0402",
  2440 => x"f4050d74",
  2441 => x"70882a83",
  2442 => x"fe800670",
  2443 => x"72982a07",
  2444 => x"72882b87",
  2445 => x"fc808006",
  2446 => x"73982b81",
  2447 => x"f00a0671",
  2448 => x"73070780",
  2449 => x"d9bc0c56",
  2450 => x"51535102",
  2451 => x"8c050d04",
  2452 => x"02f8050d",
  2453 => x"028e0580",
  2454 => x"f52d7488",
  2455 => x"2b077083",
  2456 => x"ffff0680",
  2457 => x"d9bc0c51",
  2458 => x"0288050d",
  2459 => x"0402f405",
  2460 => x"0d747678",
  2461 => x"53545280",
  2462 => x"71259738",
  2463 => x"72708105",
  2464 => x"5480f52d",
  2465 => x"72708105",
  2466 => x"5481b72d",
  2467 => x"ff115170",
  2468 => x"eb388072",
  2469 => x"81b72d02",
  2470 => x"8c050d04",
  2471 => x"02e8050d",
  2472 => x"77568070",
  2473 => x"56547376",
  2474 => x"24b73880",
  2475 => x"e1c40874",
  2476 => x"2eaf3873",
  2477 => x"5180c6e6",
  2478 => x"2d80d9bc",
  2479 => x"0880d9bc",
  2480 => x"08098105",
  2481 => x"7080d9bc",
  2482 => x"08079f2a",
  2483 => x"77058117",
  2484 => x"57575353",
  2485 => x"74762489",
  2486 => x"3880e1c4",
  2487 => x"087426d3",
  2488 => x"387280d9",
  2489 => x"bc0c0298",
  2490 => x"050d0402",
  2491 => x"f0050d80",
  2492 => x"d9b80816",
  2493 => x"5180cd9c",
  2494 => x"2d80d9bc",
  2495 => x"08802ea0",
  2496 => x"388b5380",
  2497 => x"d9bc0852",
  2498 => x"80dfb451",
  2499 => x"80cced2d",
  2500 => x"80e1f008",
  2501 => x"5473802e",
  2502 => x"873880df",
  2503 => x"b451732d",
  2504 => x"0290050d",
  2505 => x"0402dc05",
  2506 => x"0d80705a",
  2507 => x"557480d9",
  2508 => x"b80825b5",
  2509 => x"3880e1c4",
  2510 => x"08752ead",
  2511 => x"38785180",
  2512 => x"c6e62d80",
  2513 => x"d9bc0809",
  2514 => x"81057080",
  2515 => x"d9bc0807",
  2516 => x"9f2a7605",
  2517 => x"811b5b56",
  2518 => x"547480d9",
  2519 => x"b8082589",
  2520 => x"3880e1c4",
  2521 => x"087926d5",
  2522 => x"38805578",
  2523 => x"80e1c408",
  2524 => x"2781e438",
  2525 => x"785180c6",
  2526 => x"e62d80d9",
  2527 => x"bc08802e",
  2528 => x"81b43880",
  2529 => x"d9bc088b",
  2530 => x"0580f52d",
  2531 => x"70842a70",
  2532 => x"81067710",
  2533 => x"78842b80",
  2534 => x"dfb40b80",
  2535 => x"f52d5c5c",
  2536 => x"53515556",
  2537 => x"73802e80",
  2538 => x"ce387416",
  2539 => x"822b80d0",
  2540 => x"fb0b80d8",
  2541 => x"8c120c54",
  2542 => x"77753110",
  2543 => x"80e1f411",
  2544 => x"55569074",
  2545 => x"70810556",
  2546 => x"81b72da0",
  2547 => x"7481b72d",
  2548 => x"7681ff06",
  2549 => x"81165854",
  2550 => x"73802e8b",
  2551 => x"389c5380",
  2552 => x"dfb45280",
  2553 => x"cfee048b",
  2554 => x"5380d9bc",
  2555 => x"085280e1",
  2556 => x"f6165180",
  2557 => x"d0ac0474",
  2558 => x"16822b80",
  2559 => x"cdeb0b80",
  2560 => x"d88c120c",
  2561 => x"547681ff",
  2562 => x"06811658",
  2563 => x"5473802e",
  2564 => x"8b389c53",
  2565 => x"80dfb452",
  2566 => x"80d0a304",
  2567 => x"8b5380d9",
  2568 => x"bc085277",
  2569 => x"75311080",
  2570 => x"e1f40551",
  2571 => x"765580cc",
  2572 => x"ed2d80d0",
  2573 => x"cb047490",
  2574 => x"29753170",
  2575 => x"1080e1f4",
  2576 => x"05515480",
  2577 => x"d9bc0874",
  2578 => x"81b72d81",
  2579 => x"1959748b",
  2580 => x"24a43880",
  2581 => x"ceeb0474",
  2582 => x"90297531",
  2583 => x"701080e1",
  2584 => x"f4058c77",
  2585 => x"31575154",
  2586 => x"807481b7",
  2587 => x"2d9e14ff",
  2588 => x"16565474",
  2589 => x"f33802a4",
  2590 => x"050d0402",
  2591 => x"fc050d80",
  2592 => x"d9b80813",
  2593 => x"5180cd9c",
  2594 => x"2d80d9bc",
  2595 => x"08802e89",
  2596 => x"3880d9bc",
  2597 => x"0851bea5",
  2598 => x"2d800b80",
  2599 => x"d9b80c80",
  2600 => x"cea52dac",
  2601 => x"af2d0284",
  2602 => x"050d0402",
  2603 => x"fc050d72",
  2604 => x"5170fd2e",
  2605 => x"b23870fd",
  2606 => x"248b3870",
  2607 => x"fc2e80d0",
  2608 => x"3880d29a",
  2609 => x"0470fe2e",
  2610 => x"b93870ff",
  2611 => x"2e098106",
  2612 => x"80c83880",
  2613 => x"d9b80851",
  2614 => x"70802ebe",
  2615 => x"38ff1180",
  2616 => x"d9b80c80",
  2617 => x"d29a0480",
  2618 => x"d9b808f0",
  2619 => x"057080d9",
  2620 => x"b80c5170",
  2621 => x"8025a338",
  2622 => x"800b80d9",
  2623 => x"b80c80d2",
  2624 => x"9a0480d9",
  2625 => x"b8088105",
  2626 => x"80d9b80c",
  2627 => x"80d29a04",
  2628 => x"80d9b808",
  2629 => x"900580d9",
  2630 => x"b80c80ce",
  2631 => x"a52dacaf",
  2632 => x"2d028405",
  2633 => x"0d0402fc",
  2634 => x"050d800b",
  2635 => x"80d9b80c",
  2636 => x"80cea52d",
  2637 => x"abab2d80",
  2638 => x"d9bc0880",
  2639 => x"d9a80c80",
  2640 => x"d88451ad",
  2641 => x"d52d0284",
  2642 => x"050d0471",
  2643 => x"80e1f00c",
  2644 => x"04000000",
  2645 => x"00ffffff",
  2646 => x"ff00ffff",
  2647 => x"ffff00ff",
  2648 => x"ffffff00",
  2649 => x"30313233",
  2650 => x"34353637",
  2651 => x"38394142",
  2652 => x"43444546",
  2653 => x"00000000",
  2654 => x"44656275",
  2655 => x"67000000",
  2656 => x"52657365",
  2657 => x"74000000",
  2658 => x"5363616e",
  2659 => x"6c696e65",
  2660 => x"73000000",
  2661 => x"50414c20",
  2662 => x"2f204e54",
  2663 => x"53430000",
  2664 => x"436f6c6f",
  2665 => x"72000000",
  2666 => x"44696666",
  2667 => x"6963756c",
  2668 => x"74792041",
  2669 => x"00000000",
  2670 => x"44696666",
  2671 => x"6963756c",
  2672 => x"74792042",
  2673 => x"00000000",
  2674 => x"53656c65",
  2675 => x"63740000",
  2676 => x"53746172",
  2677 => x"74000000",
  2678 => x"4c6f6164",
  2679 => x"20524f4d",
  2680 => x"20100000",
  2681 => x"45786974",
  2682 => x"00000000",
  2683 => x"524f4d20",
  2684 => x"6c6f6164",
  2685 => x"696e6720",
  2686 => x"6661696c",
  2687 => x"65640000",
  2688 => x"4f4b0000",
  2689 => x"496e6974",
  2690 => x"69616c69",
  2691 => x"7a696e67",
  2692 => x"20534420",
  2693 => x"63617264",
  2694 => x"0a000000",
  2695 => x"436f6c6c",
  2696 => x"6563746f",
  2697 => x"72566973",
  2698 => x"696f6e00",
  2699 => x"16200000",
  2700 => x"14200000",
  2701 => x"15200000",
  2702 => x"53442069",
  2703 => x"6e69742e",
  2704 => x"2e2e0a00",
  2705 => x"53442063",
  2706 => x"61726420",
  2707 => x"72657365",
  2708 => x"74206661",
  2709 => x"696c6564",
  2710 => x"210a0000",
  2711 => x"53444843",
  2712 => x"20657272",
  2713 => x"6f72210a",
  2714 => x"00000000",
  2715 => x"57726974",
  2716 => x"65206661",
  2717 => x"696c6564",
  2718 => x"0a000000",
  2719 => x"52656164",
  2720 => x"20666169",
  2721 => x"6c65640a",
  2722 => x"00000000",
  2723 => x"43617264",
  2724 => x"20696e69",
  2725 => x"74206661",
  2726 => x"696c6564",
  2727 => x"0a000000",
  2728 => x"46415431",
  2729 => x"36202020",
  2730 => x"00000000",
  2731 => x"46415433",
  2732 => x"32202020",
  2733 => x"00000000",
  2734 => x"4e6f2070",
  2735 => x"61727469",
  2736 => x"74696f6e",
  2737 => x"20736967",
  2738 => x"0a000000",
  2739 => x"42616420",
  2740 => x"70617274",
  2741 => x"0a000000",
  2742 => x"4261636b",
  2743 => x"00000000",
  2744 => x"00000002",
  2745 => x"00002964",
  2746 => x"00002d28",
  2747 => x"00000002",
  2748 => x"00002ce4",
  2749 => x"000012dc",
  2750 => x"00000002",
  2751 => x"00002978",
  2752 => x"00001259",
  2753 => x"00000002",
  2754 => x"00002980",
  2755 => x"0000035a",
  2756 => x"00000001",
  2757 => x"00002988",
  2758 => x"00000000",
  2759 => x"00000001",
  2760 => x"00002994",
  2761 => x"00000001",
  2762 => x"00000001",
  2763 => x"000029a0",
  2764 => x"00000002",
  2765 => x"00000001",
  2766 => x"000029a8",
  2767 => x"00000003",
  2768 => x"00000001",
  2769 => x"000029b8",
  2770 => x"00000004",
  2771 => x"00000002",
  2772 => x"000029c8",
  2773 => x"0000036e",
  2774 => x"00000002",
  2775 => x"000029d0",
  2776 => x"00000a3f",
  2777 => x"00000002",
  2778 => x"000029d8",
  2779 => x"00002926",
  2780 => x"00000002",
  2781 => x"000029e4",
  2782 => x"000015c8",
  2783 => x"00000000",
  2784 => x"00000000",
  2785 => x"00000000",
  2786 => x"00000004",
  2787 => x"000029ec",
  2788 => x"00002b88",
  2789 => x"00000004",
  2790 => x"00002a00",
  2791 => x"00002aec",
  2792 => x"00000000",
  2793 => x"00000000",
  2794 => x"00000000",
  2795 => x"00000000",
  2796 => x"00000000",
  2797 => x"00000000",
  2798 => x"00000000",
  2799 => x"00000000",
  2800 => x"00000000",
  2801 => x"00000000",
  2802 => x"00000000",
  2803 => x"00000000",
  2804 => x"00000000",
  2805 => x"00000000",
  2806 => x"00000000",
  2807 => x"00000000",
  2808 => x"00000000",
  2809 => x"00000000",
  2810 => x"00000000",
  2811 => x"00000000",
  2812 => x"00000000",
  2813 => x"00000000",
  2814 => x"00000006",
  2815 => x"00000000",
  2816 => x"00000000",
  2817 => x"00000002",
  2818 => x"000030f4",
  2819 => x"000026eb",
  2820 => x"00000002",
  2821 => x"00003112",
  2822 => x"000026eb",
  2823 => x"00000002",
  2824 => x"00003130",
  2825 => x"000026eb",
  2826 => x"00000002",
  2827 => x"0000314e",
  2828 => x"000026eb",
  2829 => x"00000002",
  2830 => x"0000316c",
  2831 => x"000026eb",
  2832 => x"00000002",
  2833 => x"0000318a",
  2834 => x"000026eb",
  2835 => x"00000002",
  2836 => x"000031a8",
  2837 => x"000026eb",
  2838 => x"00000002",
  2839 => x"000031c6",
  2840 => x"000026eb",
  2841 => x"00000002",
  2842 => x"000031e4",
  2843 => x"000026eb",
  2844 => x"00000002",
  2845 => x"00003202",
  2846 => x"000026eb",
  2847 => x"00000002",
  2848 => x"00003220",
  2849 => x"000026eb",
  2850 => x"00000002",
  2851 => x"0000323e",
  2852 => x"000026eb",
  2853 => x"00000002",
  2854 => x"0000325c",
  2855 => x"000026eb",
  2856 => x"00000004",
  2857 => x"00002ad8",
  2858 => x"00000000",
  2859 => x"00000000",
  2860 => x"00000000",
  2861 => x"000028ab",
  2862 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

