-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80df",
     9 => x"ac080b0b",
    10 => x"80dfb008",
    11 => x"0b0b80df",
    12 => x"b4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"dfb40c0b",
    16 => x"0b80dfb0",
    17 => x"0c0b0b80",
    18 => x"dfac0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d788",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80dfac70",
    57 => x"80ebb027",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a6e1",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80df",
    65 => x"bc0c9f0b",
    66 => x"80dfc00c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"dfc008ff",
    70 => x"0580dfc0",
    71 => x"0c80dfc0",
    72 => x"088025e8",
    73 => x"3880dfbc",
    74 => x"08ff0580",
    75 => x"dfbc0c80",
    76 => x"dfbc0880",
    77 => x"25d03880",
    78 => x"0b80dfc0",
    79 => x"0c800b80",
    80 => x"dfbc0c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80dfbc08",
   100 => x"25913882",
   101 => x"c82d80df",
   102 => x"bc08ff05",
   103 => x"80dfbc0c",
   104 => x"838a0480",
   105 => x"dfbc0880",
   106 => x"dfc00853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80dfbc08",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"dfc00881",
   116 => x"0580dfc0",
   117 => x"0c80dfc0",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80dfc0",
   121 => x"0c80dfbc",
   122 => x"08810580",
   123 => x"dfbc0c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480df",
   128 => x"c0088105",
   129 => x"80dfc00c",
   130 => x"80dfc008",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80dfc0",
   134 => x"0c80dfbc",
   135 => x"08810580",
   136 => x"dfbc0c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"dfc40cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"dfc40c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280df",
   177 => x"c4088407",
   178 => x"80dfc40c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80da",
   183 => x"c40c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80dfc4",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80df",
   208 => x"ac0c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02f8050d",
  1093 => x"028f0580",
  1094 => x"f52d80da",
  1095 => x"cc085252",
  1096 => x"7080e19d",
  1097 => x"279a3871",
  1098 => x"7181b72d",
  1099 => x"80dacc08",
  1100 => x"810580da",
  1101 => x"cc0c80da",
  1102 => x"cc085180",
  1103 => x"7181b72d",
  1104 => x"0288050d",
  1105 => x"0402f405",
  1106 => x"0d747084",
  1107 => x"2a708f06",
  1108 => x"80dac808",
  1109 => x"057080f5",
  1110 => x"2d545153",
  1111 => x"53a2902d",
  1112 => x"728f0680",
  1113 => x"dac80805",
  1114 => x"7080f52d",
  1115 => x"5253a290",
  1116 => x"2d028c05",
  1117 => x"0d0402f4",
  1118 => x"050d7476",
  1119 => x"54527270",
  1120 => x"81055480",
  1121 => x"f52d5170",
  1122 => x"72708105",
  1123 => x"5481b72d",
  1124 => x"70ec3870",
  1125 => x"7281b72d",
  1126 => x"028c050d",
  1127 => x"0402d005",
  1128 => x"0d800b80",
  1129 => x"dde80881",
  1130 => x"8006715d",
  1131 => x"5d59810b",
  1132 => x"ec0c840b",
  1133 => x"ec0c7d52",
  1134 => x"80dfc851",
  1135 => x"80cdd22d",
  1136 => x"80dfac08",
  1137 => x"792e80ff",
  1138 => x"3880dfcc",
  1139 => x"0879ff12",
  1140 => x"57595774",
  1141 => x"792e8b38",
  1142 => x"81187581",
  1143 => x"2a565874",
  1144 => x"f738f718",
  1145 => x"58815980",
  1146 => x"772580db",
  1147 => x"38775274",
  1148 => x"5184a82d",
  1149 => x"80e1e852",
  1150 => x"80dfc851",
  1151 => x"80d0a82d",
  1152 => x"80dfac08",
  1153 => x"802ea638",
  1154 => x"80e1e85a",
  1155 => x"7ba73883",
  1156 => x"ff567970",
  1157 => x"81055b80",
  1158 => x"f52d7b81",
  1159 => x"1d5de40c",
  1160 => x"e80cff16",
  1161 => x"56758025",
  1162 => x"e938a4b5",
  1163 => x"0480dfac",
  1164 => x"08598480",
  1165 => x"5780dfc8",
  1166 => x"5180cff7",
  1167 => x"2dfc8017",
  1168 => x"81165657",
  1169 => x"a3e70480",
  1170 => x"dfcc08f8",
  1171 => x"0c810be0",
  1172 => x"0c805186",
  1173 => x"da2d86c7",
  1174 => x"2d78802e",
  1175 => x"883880da",
  1176 => x"d051a4e9",
  1177 => x"0480dc90",
  1178 => x"51b1f12d",
  1179 => x"7880dfac",
  1180 => x"0c02b005",
  1181 => x"0d0402ec",
  1182 => x"050d80e0",
  1183 => x"dc0b80da",
  1184 => x"cc0c80e0",
  1185 => x"dc558075",
  1186 => x"81b72d80",
  1187 => x"dcb40851",
  1188 => x"a2c52dba",
  1189 => x"51a2902d",
  1190 => x"ffb408ff",
  1191 => x"b8087098",
  1192 => x"2a535154",
  1193 => x"a2c52d73",
  1194 => x"902a7081",
  1195 => x"ff065253",
  1196 => x"a2c52d73",
  1197 => x"882a7081",
  1198 => x"ff065253",
  1199 => x"a2c52d73",
  1200 => x"81ff0651",
  1201 => x"a2c52d74",
  1202 => x"5280dfd4",
  1203 => x"51a2f62d",
  1204 => x"7480dacc",
  1205 => x"0c807581",
  1206 => x"b72d80dd",
  1207 => x"8c707070",
  1208 => x"84055208",
  1209 => x"535454a2",
  1210 => x"c52d7208",
  1211 => x"51a2c52d",
  1212 => x"88140851",
  1213 => x"a2c52d80",
  1214 => x"dacc0853",
  1215 => x"a07381b7",
  1216 => x"2d80dacc",
  1217 => x"08810580",
  1218 => x"dacc0c8c",
  1219 => x"140851a2",
  1220 => x"c52d9014",
  1221 => x"0851a2c5",
  1222 => x"2d941408",
  1223 => x"51a2c52d",
  1224 => x"80dacc08",
  1225 => x"53a07381",
  1226 => x"b72d80da",
  1227 => x"cc088105",
  1228 => x"80dacc0c",
  1229 => x"98140851",
  1230 => x"a2c52d74",
  1231 => x"5280e098",
  1232 => x"51a2f62d",
  1233 => x"80dad051",
  1234 => x"b1f12d80",
  1235 => x"dcb40884",
  1236 => x"0580dcb4",
  1237 => x"0c029405",
  1238 => x"0d04800b",
  1239 => x"80dcb40c",
  1240 => x"0402ec05",
  1241 => x"0d840bec",
  1242 => x"0cafae2d",
  1243 => x"a9972d81",
  1244 => x"f92d8353",
  1245 => x"af912d81",
  1246 => x"51858d2d",
  1247 => x"ff135372",
  1248 => x"8025f138",
  1249 => x"840bec0c",
  1250 => x"80d8e051",
  1251 => x"86a02d80",
  1252 => x"c3f32d80",
  1253 => x"dfac0880",
  1254 => x"2e81e538",
  1255 => x"a39d5180",
  1256 => x"d6ff2d80",
  1257 => x"d8f85280",
  1258 => x"dfd451a2",
  1259 => x"f62d80d9",
  1260 => x"885280e0",
  1261 => x"9851a2f6",
  1262 => x"2d80dad0",
  1263 => x"51b1f12d",
  1264 => x"afd02daa",
  1265 => x"c22d80df",
  1266 => x"ac088106",
  1267 => x"5372802e",
  1268 => x"86388051",
  1269 => x"94bf2db2",
  1270 => x"842d80da",
  1271 => x"e40b80f5",
  1272 => x"2d80dde8",
  1273 => x"08708106",
  1274 => x"55565472",
  1275 => x"802e8538",
  1276 => x"73840754",
  1277 => x"74812a70",
  1278 => x"81065153",
  1279 => x"72802e85",
  1280 => x"38738207",
  1281 => x"5474822a",
  1282 => x"70810651",
  1283 => x"5372802e",
  1284 => x"85387381",
  1285 => x"07547483",
  1286 => x"2a708106",
  1287 => x"51537280",
  1288 => x"2e853873",
  1289 => x"88075474",
  1290 => x"842a7081",
  1291 => x"06515372",
  1292 => x"802e8538",
  1293 => x"73900754",
  1294 => x"74852a70",
  1295 => x"81065153",
  1296 => x"72802e85",
  1297 => x"3873a007",
  1298 => x"5474882a",
  1299 => x"70810651",
  1300 => x"5372802e",
  1301 => x"86387380",
  1302 => x"c0075474",
  1303 => x"892a7081",
  1304 => x"06515372",
  1305 => x"802e8638",
  1306 => x"73818007",
  1307 => x"5473fc0c",
  1308 => x"865380df",
  1309 => x"ac088338",
  1310 => x"845372ec",
  1311 => x"0ca7c304",
  1312 => x"800b80df",
  1313 => x"ac0c0294",
  1314 => x"050d0471",
  1315 => x"980c04ff",
  1316 => x"b00880df",
  1317 => x"ac0c0481",
  1318 => x"0bffb00c",
  1319 => x"04800bff",
  1320 => x"b00c0402",
  1321 => x"d8050dff",
  1322 => x"b40887ff",
  1323 => x"ff065a81",
  1324 => x"54807080",
  1325 => x"ddd40880",
  1326 => x"ddd80880",
  1327 => x"ddb05b59",
  1328 => x"575a5879",
  1329 => x"74067575",
  1330 => x"06525271",
  1331 => x"712e8d38",
  1332 => x"8077818a",
  1333 => x"2d730975",
  1334 => x"06720755",
  1335 => x"7680e02d",
  1336 => x"7083ffff",
  1337 => x"06535171",
  1338 => x"83f42e09",
  1339 => x"8106a238",
  1340 => x"74740670",
  1341 => x"77760632",
  1342 => x"70098105",
  1343 => x"7072079f",
  1344 => x"2a7b0577",
  1345 => x"097a0674",
  1346 => x"075a5b53",
  1347 => x"5353aa9f",
  1348 => x"047183f4",
  1349 => x"26893881",
  1350 => x"11517077",
  1351 => x"818a2d73",
  1352 => x"10811a82",
  1353 => x"19595a54",
  1354 => x"907925ff",
  1355 => x"96387580",
  1356 => x"ddd80c74",
  1357 => x"80ddd40c",
  1358 => x"7780dfac",
  1359 => x"0c02a805",
  1360 => x"0d0402cc",
  1361 => x"050d805d",
  1362 => x"abd20480",
  1363 => x"dfac0881",
  1364 => x"f02e0981",
  1365 => x"068a3881",
  1366 => x"0b80dde0",
  1367 => x"0cabd204",
  1368 => x"80dfac08",
  1369 => x"81e02e09",
  1370 => x"81068a38",
  1371 => x"810b80dd",
  1372 => x"e40cabd2",
  1373 => x"0480dfac",
  1374 => x"085280dd",
  1375 => x"e408802e",
  1376 => x"893880df",
  1377 => x"ac088180",
  1378 => x"05527184",
  1379 => x"2c728f06",
  1380 => x"535380dd",
  1381 => x"e008802e",
  1382 => x"9a387284",
  1383 => x"2980dcb8",
  1384 => x"05721381",
  1385 => x"712b7009",
  1386 => x"73080673",
  1387 => x"0c515353",
  1388 => x"abc60472",
  1389 => x"842980dc",
  1390 => x"b8057213",
  1391 => x"83712b72",
  1392 => x"0807720c",
  1393 => x"5353800b",
  1394 => x"80dde40c",
  1395 => x"800b80dd",
  1396 => x"e00c80e1",
  1397 => x"a051ae84",
  1398 => x"2d80dfac",
  1399 => x"08ff24fe",
  1400 => x"ea38a9a3",
  1401 => x"2d80dfac",
  1402 => x"08802e81",
  1403 => x"a138815a",
  1404 => x"800b80dd",
  1405 => x"dc0880dd",
  1406 => x"d80880dd",
  1407 => x"e00880dd",
  1408 => x"8c5c5a5d",
  1409 => x"5d597b7a",
  1410 => x"067b7b06",
  1411 => x"57527176",
  1412 => x"2e80df38",
  1413 => x"7580dcf8",
  1414 => x"1a80f52d",
  1415 => x"70842c71",
  1416 => x"8f065754",
  1417 => x"56577580",
  1418 => x"2ea63871",
  1419 => x"842980dc",
  1420 => x"b8057415",
  1421 => x"81712b70",
  1422 => x"09730806",
  1423 => x"730c5154",
  1424 => x"527780e0",
  1425 => x"2d810552",
  1426 => x"7178818a",
  1427 => x"2dace304",
  1428 => x"71842980",
  1429 => x"dcb80574",
  1430 => x"1583712b",
  1431 => x"72080772",
  1432 => x"0c535374",
  1433 => x"852e0981",
  1434 => x"06883875",
  1435 => x"802e8338",
  1436 => x"815d7910",
  1437 => x"811a821a",
  1438 => x"5a5a5a90",
  1439 => x"7925ff86",
  1440 => x"387680dd",
  1441 => x"e00c80dd",
  1442 => x"d80880dd",
  1443 => x"dc0c7c80",
  1444 => x"dfac0c02",
  1445 => x"b4050d04",
  1446 => x"02f8050d",
  1447 => x"80dcb852",
  1448 => x"8f518072",
  1449 => x"70840554",
  1450 => x"0cff1151",
  1451 => x"708025f2",
  1452 => x"38028805",
  1453 => x"0d0402f0",
  1454 => x"050d7551",
  1455 => x"a99d2d70",
  1456 => x"822cfc06",
  1457 => x"80dcb811",
  1458 => x"72109e06",
  1459 => x"71087072",
  1460 => x"2a708306",
  1461 => x"82742b70",
  1462 => x"09740676",
  1463 => x"0c545156",
  1464 => x"57535153",
  1465 => x"a9972d71",
  1466 => x"80dfac0c",
  1467 => x"0290050d",
  1468 => x"0402fc05",
  1469 => x"0d725180",
  1470 => x"710c800b",
  1471 => x"84120c02",
  1472 => x"84050d04",
  1473 => x"02f0050d",
  1474 => x"75700884",
  1475 => x"12085353",
  1476 => x"53ff5471",
  1477 => x"712ea838",
  1478 => x"a99d2d84",
  1479 => x"13087084",
  1480 => x"29148811",
  1481 => x"70087081",
  1482 => x"ff068418",
  1483 => x"08811187",
  1484 => x"06841a0c",
  1485 => x"53515551",
  1486 => x"5151a997",
  1487 => x"2d715473",
  1488 => x"80dfac0c",
  1489 => x"0290050d",
  1490 => x"0402f805",
  1491 => x"0da99d2d",
  1492 => x"e008708b",
  1493 => x"2a708106",
  1494 => x"51525270",
  1495 => x"802ea138",
  1496 => x"80e1a008",
  1497 => x"70842980",
  1498 => x"e1a80573",
  1499 => x"81ff0671",
  1500 => x"0c515180",
  1501 => x"e1a00881",
  1502 => x"11870680",
  1503 => x"e1a00c51",
  1504 => x"800b80e1",
  1505 => x"c80ca98f",
  1506 => x"2da9972d",
  1507 => x"0288050d",
  1508 => x"0402fc05",
  1509 => x"0da99d2d",
  1510 => x"810b80e1",
  1511 => x"c80ca997",
  1512 => x"2d80e1c8",
  1513 => x"085170f9",
  1514 => x"38028405",
  1515 => x"0d0402fc",
  1516 => x"050d80e1",
  1517 => x"a051adf1",
  1518 => x"2dad982d",
  1519 => x"aec951a9",
  1520 => x"8b2d0284",
  1521 => x"050d0480",
  1522 => x"e1d40880",
  1523 => x"dfac0c04",
  1524 => x"02fc050d",
  1525 => x"810b80dd",
  1526 => x"ec0c8151",
  1527 => x"858d2d02",
  1528 => x"84050d04",
  1529 => x"02fc050d",
  1530 => x"afee04aa",
  1531 => x"c22d80f6",
  1532 => x"51adb62d",
  1533 => x"80dfac08",
  1534 => x"f23880da",
  1535 => x"51adb62d",
  1536 => x"80dfac08",
  1537 => x"e63880df",
  1538 => x"ac0880dd",
  1539 => x"ec0c80df",
  1540 => x"ac085185",
  1541 => x"8d2d0284",
  1542 => x"050d0402",
  1543 => x"ec050d76",
  1544 => x"54805287",
  1545 => x"0b881580",
  1546 => x"f52d5653",
  1547 => x"74722483",
  1548 => x"38a05372",
  1549 => x"5183842d",
  1550 => x"81128b15",
  1551 => x"80f52d54",
  1552 => x"52727225",
  1553 => x"de380294",
  1554 => x"050d0402",
  1555 => x"f0050d80",
  1556 => x"e1d40854",
  1557 => x"81f92d80",
  1558 => x"0b80e1d8",
  1559 => x"0c730880",
  1560 => x"2e818938",
  1561 => x"820b80df",
  1562 => x"c00c80e1",
  1563 => x"d8088f06",
  1564 => x"80dfbc0c",
  1565 => x"73085271",
  1566 => x"832e9638",
  1567 => x"71832689",
  1568 => x"3871812e",
  1569 => x"b038b1d5",
  1570 => x"0471852e",
  1571 => x"a038b1d5",
  1572 => x"04881480",
  1573 => x"f52d8415",
  1574 => x"0880d990",
  1575 => x"53545286",
  1576 => x"a02d7184",
  1577 => x"29137008",
  1578 => x"5252b1d9",
  1579 => x"047351b0",
  1580 => x"9b2db1d5",
  1581 => x"0480dde8",
  1582 => x"08881508",
  1583 => x"2c708106",
  1584 => x"51527180",
  1585 => x"2e883880",
  1586 => x"d99451b1",
  1587 => x"d20480d9",
  1588 => x"985186a0",
  1589 => x"2d841408",
  1590 => x"5186a02d",
  1591 => x"80e1d808",
  1592 => x"810580e1",
  1593 => x"d80c8c14",
  1594 => x"54b0dd04",
  1595 => x"0290050d",
  1596 => x"047180e1",
  1597 => x"d40cb0cb",
  1598 => x"2d80e1d8",
  1599 => x"08ff0580",
  1600 => x"e1dc0c04",
  1601 => x"02e8050d",
  1602 => x"80e1d408",
  1603 => x"80e1e008",
  1604 => x"575580f6",
  1605 => x"51adb62d",
  1606 => x"80dfac08",
  1607 => x"812a7081",
  1608 => x"06515271",
  1609 => x"802ea438",
  1610 => x"b2ae04aa",
  1611 => x"c22d80f6",
  1612 => x"51adb62d",
  1613 => x"80dfac08",
  1614 => x"f23880dd",
  1615 => x"ec088132",
  1616 => x"7080ddec",
  1617 => x"0c705252",
  1618 => x"858d2d80",
  1619 => x"0b80e1cc",
  1620 => x"0c800b80",
  1621 => x"e1d00c80",
  1622 => x"ddec0883",
  1623 => x"8d3880da",
  1624 => x"51adb62d",
  1625 => x"80dfac08",
  1626 => x"802e8c38",
  1627 => x"80e1cc08",
  1628 => x"81800780",
  1629 => x"e1cc0c80",
  1630 => x"d951adb6",
  1631 => x"2d80dfac",
  1632 => x"08802e8c",
  1633 => x"3880e1cc",
  1634 => x"0880c007",
  1635 => x"80e1cc0c",
  1636 => x"819451ad",
  1637 => x"b62d80df",
  1638 => x"ac08802e",
  1639 => x"8b3880e1",
  1640 => x"cc089007",
  1641 => x"80e1cc0c",
  1642 => x"819151ad",
  1643 => x"b62d80df",
  1644 => x"ac08802e",
  1645 => x"8b3880e1",
  1646 => x"cc08a007",
  1647 => x"80e1cc0c",
  1648 => x"81f551ad",
  1649 => x"b62d80df",
  1650 => x"ac08802e",
  1651 => x"8b3880e1",
  1652 => x"cc088107",
  1653 => x"80e1cc0c",
  1654 => x"81f251ad",
  1655 => x"b62d80df",
  1656 => x"ac08802e",
  1657 => x"8b3880e1",
  1658 => x"cc088207",
  1659 => x"80e1cc0c",
  1660 => x"81eb51ad",
  1661 => x"b62d80df",
  1662 => x"ac08802e",
  1663 => x"8b3880e1",
  1664 => x"cc088407",
  1665 => x"80e1cc0c",
  1666 => x"81f451ad",
  1667 => x"b62d80df",
  1668 => x"ac08802e",
  1669 => x"8b3880e1",
  1670 => x"cc088807",
  1671 => x"80e1cc0c",
  1672 => x"80d851ad",
  1673 => x"b62d80df",
  1674 => x"ac08802e",
  1675 => x"8c3880e1",
  1676 => x"d0088180",
  1677 => x"0780e1d0",
  1678 => x"0c9251ad",
  1679 => x"b62d80df",
  1680 => x"ac08802e",
  1681 => x"8c3880e1",
  1682 => x"d00880c0",
  1683 => x"0780e1d0",
  1684 => x"0c9451ad",
  1685 => x"b62d80df",
  1686 => x"ac08802e",
  1687 => x"8b3880e1",
  1688 => x"d0089007",
  1689 => x"80e1d00c",
  1690 => x"9151adb6",
  1691 => x"2d80dfac",
  1692 => x"08802e8b",
  1693 => x"3880e1d0",
  1694 => x"08a00780",
  1695 => x"e1d00c9d",
  1696 => x"51adb62d",
  1697 => x"80dfac08",
  1698 => x"802e8b38",
  1699 => x"80e1d008",
  1700 => x"810780e1",
  1701 => x"d00c9b51",
  1702 => x"adb62d80",
  1703 => x"dfac0880",
  1704 => x"2e8b3880",
  1705 => x"e1d00882",
  1706 => x"0780e1d0",
  1707 => x"0c9c51ad",
  1708 => x"b62d80df",
  1709 => x"ac08802e",
  1710 => x"8b3880e1",
  1711 => x"d0088407",
  1712 => x"80e1d00c",
  1713 => x"a351adb6",
  1714 => x"2d80dfac",
  1715 => x"08802e8b",
  1716 => x"3880e1d0",
  1717 => x"08880780",
  1718 => x"e1d00c81",
  1719 => x"fd51adb6",
  1720 => x"2d81fa51",
  1721 => x"adb62dbb",
  1722 => x"bf0481f5",
  1723 => x"51adb62d",
  1724 => x"80dfac08",
  1725 => x"812a7081",
  1726 => x"06515271",
  1727 => x"802eb338",
  1728 => x"80e1dc08",
  1729 => x"5271802e",
  1730 => x"8a38ff12",
  1731 => x"80e1dc0c",
  1732 => x"b6b20480",
  1733 => x"e1d80810",
  1734 => x"80e1d808",
  1735 => x"05708429",
  1736 => x"16515288",
  1737 => x"1208802e",
  1738 => x"8938ff51",
  1739 => x"88120852",
  1740 => x"712d81f2",
  1741 => x"51adb62d",
  1742 => x"80dfac08",
  1743 => x"812a7081",
  1744 => x"06515271",
  1745 => x"802eb438",
  1746 => x"80e1d808",
  1747 => x"ff1180e1",
  1748 => x"dc085653",
  1749 => x"53737225",
  1750 => x"8a388114",
  1751 => x"80e1dc0c",
  1752 => x"b6fb0472",
  1753 => x"10137084",
  1754 => x"29165152",
  1755 => x"88120880",
  1756 => x"2e8938fe",
  1757 => x"51881208",
  1758 => x"52712d81",
  1759 => x"fd51adb6",
  1760 => x"2d80dfac",
  1761 => x"08812a70",
  1762 => x"81065152",
  1763 => x"71802eb1",
  1764 => x"3880e1dc",
  1765 => x"08802e8a",
  1766 => x"38800b80",
  1767 => x"e1dc0cb7",
  1768 => x"c10480e1",
  1769 => x"d8081080",
  1770 => x"e1d80805",
  1771 => x"70842916",
  1772 => x"51528812",
  1773 => x"08802e89",
  1774 => x"38fd5188",
  1775 => x"12085271",
  1776 => x"2d81fa51",
  1777 => x"adb62d80",
  1778 => x"dfac0881",
  1779 => x"2a708106",
  1780 => x"51527180",
  1781 => x"2eb13880",
  1782 => x"e1d808ff",
  1783 => x"11545280",
  1784 => x"e1dc0873",
  1785 => x"25893872",
  1786 => x"80e1dc0c",
  1787 => x"b8870471",
  1788 => x"10127084",
  1789 => x"29165152",
  1790 => x"88120880",
  1791 => x"2e8938fc",
  1792 => x"51881208",
  1793 => x"52712d80",
  1794 => x"e1dc0870",
  1795 => x"53547380",
  1796 => x"2e8a388c",
  1797 => x"15ff1555",
  1798 => x"55b88e04",
  1799 => x"820b80df",
  1800 => x"c00c718f",
  1801 => x"0680dfbc",
  1802 => x"0c81eb51",
  1803 => x"adb62d80",
  1804 => x"dfac0881",
  1805 => x"2a708106",
  1806 => x"51527180",
  1807 => x"2ead3874",
  1808 => x"08852e09",
  1809 => x"8106a438",
  1810 => x"881580f5",
  1811 => x"2dff0552",
  1812 => x"71881681",
  1813 => x"b72d7198",
  1814 => x"2b527180",
  1815 => x"25883880",
  1816 => x"0b881681",
  1817 => x"b72d7451",
  1818 => x"b09b2d81",
  1819 => x"f451adb6",
  1820 => x"2d80dfac",
  1821 => x"08812a70",
  1822 => x"81065152",
  1823 => x"71802eb3",
  1824 => x"38740885",
  1825 => x"2e098106",
  1826 => x"aa388815",
  1827 => x"80f52d81",
  1828 => x"05527188",
  1829 => x"1681b72d",
  1830 => x"7181ff06",
  1831 => x"8b1680f5",
  1832 => x"2d545272",
  1833 => x"72278738",
  1834 => x"72881681",
  1835 => x"b72d7451",
  1836 => x"b09b2d80",
  1837 => x"da51adb6",
  1838 => x"2d80dfac",
  1839 => x"08812a70",
  1840 => x"81065152",
  1841 => x"71802e81",
  1842 => x"ad3880e1",
  1843 => x"d40880e1",
  1844 => x"dc085553",
  1845 => x"73802e8a",
  1846 => x"388c13ff",
  1847 => x"155553b9",
  1848 => x"d4047208",
  1849 => x"5271822e",
  1850 => x"a6387182",
  1851 => x"26893871",
  1852 => x"812eaa38",
  1853 => x"baf60471",
  1854 => x"832eb438",
  1855 => x"71842e09",
  1856 => x"810680f2",
  1857 => x"38881308",
  1858 => x"51b1f12d",
  1859 => x"baf60480",
  1860 => x"e1dc0851",
  1861 => x"88130852",
  1862 => x"712dbaf6",
  1863 => x"04810b88",
  1864 => x"14082b80",
  1865 => x"dde80832",
  1866 => x"80dde80c",
  1867 => x"baca0488",
  1868 => x"1380f52d",
  1869 => x"81058b14",
  1870 => x"80f52d53",
  1871 => x"54717424",
  1872 => x"83388054",
  1873 => x"73881481",
  1874 => x"b72db0cb",
  1875 => x"2dbaf604",
  1876 => x"7508802e",
  1877 => x"a4387508",
  1878 => x"51adb62d",
  1879 => x"80dfac08",
  1880 => x"81065271",
  1881 => x"802e8c38",
  1882 => x"80e1dc08",
  1883 => x"51841608",
  1884 => x"52712d88",
  1885 => x"165675d8",
  1886 => x"38805480",
  1887 => x"0b80dfc0",
  1888 => x"0c738f06",
  1889 => x"80dfbc0c",
  1890 => x"a0527380",
  1891 => x"e1dc082e",
  1892 => x"09810699",
  1893 => x"3880e1d8",
  1894 => x"08ff0574",
  1895 => x"32700981",
  1896 => x"05707207",
  1897 => x"9f2a9171",
  1898 => x"31515153",
  1899 => x"53715183",
  1900 => x"842d8114",
  1901 => x"548e7425",
  1902 => x"c23880dd",
  1903 => x"ec085271",
  1904 => x"80dfac0c",
  1905 => x"0298050d",
  1906 => x"0402f405",
  1907 => x"0dd45281",
  1908 => x"ff720c71",
  1909 => x"085381ff",
  1910 => x"720c7288",
  1911 => x"2b83fe80",
  1912 => x"06720870",
  1913 => x"81ff0651",
  1914 => x"525381ff",
  1915 => x"720c7271",
  1916 => x"07882b72",
  1917 => x"087081ff",
  1918 => x"06515253",
  1919 => x"81ff720c",
  1920 => x"72710788",
  1921 => x"2b720870",
  1922 => x"81ff0672",
  1923 => x"0780dfac",
  1924 => x"0c525302",
  1925 => x"8c050d04",
  1926 => x"02f4050d",
  1927 => x"74767181",
  1928 => x"ff06d40c",
  1929 => x"535380e1",
  1930 => x"e4088538",
  1931 => x"71892b52",
  1932 => x"71982ad4",
  1933 => x"0c71902a",
  1934 => x"7081ff06",
  1935 => x"d40c5171",
  1936 => x"882a7081",
  1937 => x"ff06d40c",
  1938 => x"517181ff",
  1939 => x"06d40c72",
  1940 => x"902a7081",
  1941 => x"ff06d40c",
  1942 => x"51d40870",
  1943 => x"81ff0651",
  1944 => x"5182b8bf",
  1945 => x"527081ff",
  1946 => x"2e098106",
  1947 => x"943881ff",
  1948 => x"0bd40cd4",
  1949 => x"087081ff",
  1950 => x"06ff1454",
  1951 => x"515171e5",
  1952 => x"387080df",
  1953 => x"ac0c028c",
  1954 => x"050d0402",
  1955 => x"fc050d81",
  1956 => x"c75181ff",
  1957 => x"0bd40cff",
  1958 => x"11517080",
  1959 => x"25f43802",
  1960 => x"84050d04",
  1961 => x"02f4050d",
  1962 => x"81ff0bd4",
  1963 => x"0c935380",
  1964 => x"5287fc80",
  1965 => x"c151bc98",
  1966 => x"2d80dfac",
  1967 => x"088b3881",
  1968 => x"ff0bd40c",
  1969 => x"8153bdd2",
  1970 => x"04bd8b2d",
  1971 => x"ff135372",
  1972 => x"de387280",
  1973 => x"dfac0c02",
  1974 => x"8c050d04",
  1975 => x"02ec050d",
  1976 => x"810b80e1",
  1977 => x"e40c8454",
  1978 => x"d008708f",
  1979 => x"2a708106",
  1980 => x"51515372",
  1981 => x"f33872d0",
  1982 => x"0cbd8b2d",
  1983 => x"80d99c51",
  1984 => x"86a02dd0",
  1985 => x"08708f2a",
  1986 => x"70810651",
  1987 => x"515372f3",
  1988 => x"38810bd0",
  1989 => x"0cb15380",
  1990 => x"5284d480",
  1991 => x"c051bc98",
  1992 => x"2d80dfac",
  1993 => x"08812e93",
  1994 => x"3872822e",
  1995 => x"bf38ff13",
  1996 => x"5372e438",
  1997 => x"ff145473",
  1998 => x"ffae38bd",
  1999 => x"8b2d83aa",
  2000 => x"52849c80",
  2001 => x"c851bc98",
  2002 => x"2d80dfac",
  2003 => x"08812e09",
  2004 => x"81069338",
  2005 => x"bbc92d80",
  2006 => x"dfac0883",
  2007 => x"ffff0653",
  2008 => x"7283aa2e",
  2009 => x"a138bda4",
  2010 => x"2dbf8004",
  2011 => x"80d9a851",
  2012 => x"86a02d80",
  2013 => x"5380c0d8",
  2014 => x"0480d9c0",
  2015 => x"5186a02d",
  2016 => x"805480c0",
  2017 => x"a90481ff",
  2018 => x"0bd40cb1",
  2019 => x"54bd8b2d",
  2020 => x"8fcf5380",
  2021 => x"5287fc80",
  2022 => x"f751bc98",
  2023 => x"2d80dfac",
  2024 => x"085580df",
  2025 => x"ac08812e",
  2026 => x"0981069c",
  2027 => x"3881ff0b",
  2028 => x"d40c820a",
  2029 => x"52849c80",
  2030 => x"e951bc98",
  2031 => x"2d80dfac",
  2032 => x"08802e8e",
  2033 => x"38bd8b2d",
  2034 => x"ff135372",
  2035 => x"c63880c0",
  2036 => x"9c0481ff",
  2037 => x"0bd40c80",
  2038 => x"dfac0852",
  2039 => x"87fc80fa",
  2040 => x"51bc982d",
  2041 => x"80dfac08",
  2042 => x"b33881ff",
  2043 => x"0bd40cd4",
  2044 => x"085381ff",
  2045 => x"0bd40c81",
  2046 => x"ff0bd40c",
  2047 => x"81ff0bd4",
  2048 => x"0c81ff0b",
  2049 => x"d40c7286",
  2050 => x"2a708106",
  2051 => x"76565153",
  2052 => x"72973880",
  2053 => x"dfac0854",
  2054 => x"80c0a904",
  2055 => x"73822efe",
  2056 => x"d838ff14",
  2057 => x"5473fee5",
  2058 => x"387380e1",
  2059 => x"e40c738b",
  2060 => x"38815287",
  2061 => x"fc80d051",
  2062 => x"bc982d81",
  2063 => x"ff0bd40c",
  2064 => x"d008708f",
  2065 => x"2a708106",
  2066 => x"51515372",
  2067 => x"f33872d0",
  2068 => x"0c81ff0b",
  2069 => x"d40c8153",
  2070 => x"7280dfac",
  2071 => x"0c029405",
  2072 => x"0d0402e8",
  2073 => x"050d7855",
  2074 => x"805681ff",
  2075 => x"0bd40cd0",
  2076 => x"08708f2a",
  2077 => x"70810651",
  2078 => x"515372f3",
  2079 => x"3882810b",
  2080 => x"d00c81ff",
  2081 => x"0bd40c77",
  2082 => x"5287fc80",
  2083 => x"d151bc98",
  2084 => x"2d80dbc6",
  2085 => x"df5480df",
  2086 => x"ac08802e",
  2087 => x"8c3880d9",
  2088 => x"e05186a0",
  2089 => x"2d80c1fe",
  2090 => x"0481ff0b",
  2091 => x"d40cd408",
  2092 => x"7081ff06",
  2093 => x"51537281",
  2094 => x"fe2e0981",
  2095 => x"069f3880",
  2096 => x"ff53bbc9",
  2097 => x"2d80dfac",
  2098 => x"08757084",
  2099 => x"05570cff",
  2100 => x"13537280",
  2101 => x"25ec3881",
  2102 => x"5680c1e3",
  2103 => x"04ff1454",
  2104 => x"73c73881",
  2105 => x"ff0bd40c",
  2106 => x"81ff0bd4",
  2107 => x"0cd00870",
  2108 => x"8f2a7081",
  2109 => x"06515153",
  2110 => x"72f33872",
  2111 => x"d00c7580",
  2112 => x"dfac0c02",
  2113 => x"98050d04",
  2114 => x"02e8050d",
  2115 => x"77797b58",
  2116 => x"55558053",
  2117 => x"727625a5",
  2118 => x"38747081",
  2119 => x"055680f5",
  2120 => x"2d747081",
  2121 => x"055680f5",
  2122 => x"2d525271",
  2123 => x"712e8738",
  2124 => x"815180c2",
  2125 => x"bf048113",
  2126 => x"5380c294",
  2127 => x"04805170",
  2128 => x"80dfac0c",
  2129 => x"0298050d",
  2130 => x"0402ec05",
  2131 => x"0d765574",
  2132 => x"802e80c4",
  2133 => x"389a1580",
  2134 => x"e02d5180",
  2135 => x"d1832d80",
  2136 => x"dfac0880",
  2137 => x"dfac0880",
  2138 => x"e8980c80",
  2139 => x"dfac0854",
  2140 => x"5480e7f4",
  2141 => x"08802e9b",
  2142 => x"38941580",
  2143 => x"e02d5180",
  2144 => x"d1832d80",
  2145 => x"dfac0890",
  2146 => x"2b83fff0",
  2147 => x"0a067075",
  2148 => x"07515372",
  2149 => x"80e8980c",
  2150 => x"80e89808",
  2151 => x"5372802e",
  2152 => x"9e3880e7",
  2153 => x"ec08fe14",
  2154 => x"712980e8",
  2155 => x"80080580",
  2156 => x"e89c0c70",
  2157 => x"842b80e7",
  2158 => x"f80c5480",
  2159 => x"c3ee0480",
  2160 => x"e8840880",
  2161 => x"e8980c80",
  2162 => x"e8880880",
  2163 => x"e89c0c80",
  2164 => x"e7f40880",
  2165 => x"2e8c3880",
  2166 => x"e7ec0884",
  2167 => x"2b5380c3",
  2168 => x"e90480e8",
  2169 => x"8c08842b",
  2170 => x"537280e7",
  2171 => x"f80c0294",
  2172 => x"050d0402",
  2173 => x"d8050d80",
  2174 => x"0b80e7f4",
  2175 => x"0c8454bd",
  2176 => x"dc2d80df",
  2177 => x"ac08802e",
  2178 => x"993880e1",
  2179 => x"e8528051",
  2180 => x"80c0e22d",
  2181 => x"80dfac08",
  2182 => x"802e8738",
  2183 => x"fe5480c4",
  2184 => x"aa04ff14",
  2185 => x"54738024",
  2186 => x"d638738e",
  2187 => x"3880d9f0",
  2188 => x"5186a02d",
  2189 => x"735580ca",
  2190 => x"8e048056",
  2191 => x"810b80e8",
  2192 => x"a00c8853",
  2193 => x"80da8452",
  2194 => x"80e29e51",
  2195 => x"80c2882d",
  2196 => x"80dfac08",
  2197 => x"762e0981",
  2198 => x"06893880",
  2199 => x"dfac0880",
  2200 => x"e8a00c88",
  2201 => x"5380da90",
  2202 => x"5280e2ba",
  2203 => x"5180c288",
  2204 => x"2d80dfac",
  2205 => x"08893880",
  2206 => x"dfac0880",
  2207 => x"e8a00c80",
  2208 => x"e8a00880",
  2209 => x"2e818538",
  2210 => x"80e5ae0b",
  2211 => x"80f52d80",
  2212 => x"e5af0b80",
  2213 => x"f52d7198",
  2214 => x"2b71902b",
  2215 => x"0780e5b0",
  2216 => x"0b80f52d",
  2217 => x"70882b72",
  2218 => x"0780e5b1",
  2219 => x"0b80f52d",
  2220 => x"710780e5",
  2221 => x"e60b80f5",
  2222 => x"2d80e5e7",
  2223 => x"0b80f52d",
  2224 => x"71882b07",
  2225 => x"535f5452",
  2226 => x"5a565755",
  2227 => x"7381abaa",
  2228 => x"2e098106",
  2229 => x"90387551",
  2230 => x"80d0d22d",
  2231 => x"80dfac08",
  2232 => x"5680c5f4",
  2233 => x"047382d4",
  2234 => x"d52e8938",
  2235 => x"80da9c51",
  2236 => x"80c6c404",
  2237 => x"80e1e852",
  2238 => x"755180c0",
  2239 => x"e22d80df",
  2240 => x"ac085580",
  2241 => x"dfac0880",
  2242 => x"2e848338",
  2243 => x"885380da",
  2244 => x"905280e2",
  2245 => x"ba5180c2",
  2246 => x"882d80df",
  2247 => x"ac088b38",
  2248 => x"810b80e7",
  2249 => x"f40c80c6",
  2250 => x"cb048853",
  2251 => x"80da8452",
  2252 => x"80e29e51",
  2253 => x"80c2882d",
  2254 => x"80dfac08",
  2255 => x"802e8c38",
  2256 => x"80dab051",
  2257 => x"86a02d80",
  2258 => x"c7aa0480",
  2259 => x"e5e60b80",
  2260 => x"f52d5473",
  2261 => x"80d52e09",
  2262 => x"810680ce",
  2263 => x"3880e5e7",
  2264 => x"0b80f52d",
  2265 => x"547381aa",
  2266 => x"2e098106",
  2267 => x"bd38800b",
  2268 => x"80e1e80b",
  2269 => x"80f52d56",
  2270 => x"547481e9",
  2271 => x"2e833881",
  2272 => x"547481eb",
  2273 => x"2e8c3880",
  2274 => x"5573752e",
  2275 => x"09810682",
  2276 => x"fd3880e1",
  2277 => x"f30b80f5",
  2278 => x"2d55748e",
  2279 => x"3880e1f4",
  2280 => x"0b80f52d",
  2281 => x"5473822e",
  2282 => x"87388055",
  2283 => x"80ca8e04",
  2284 => x"80e1f50b",
  2285 => x"80f52d70",
  2286 => x"80e7ec0c",
  2287 => x"ff0580e7",
  2288 => x"f00c80e1",
  2289 => x"f60b80f5",
  2290 => x"2d80e1f7",
  2291 => x"0b80f52d",
  2292 => x"58760577",
  2293 => x"82802905",
  2294 => x"7080e7fc",
  2295 => x"0c80e1f8",
  2296 => x"0b80f52d",
  2297 => x"7080e890",
  2298 => x"0c80e7f4",
  2299 => x"08595758",
  2300 => x"76802e81",
  2301 => x"b9388853",
  2302 => x"80da9052",
  2303 => x"80e2ba51",
  2304 => x"80c2882d",
  2305 => x"80dfac08",
  2306 => x"82843880",
  2307 => x"e7ec0870",
  2308 => x"842b80e7",
  2309 => x"f80c7080",
  2310 => x"e88c0c80",
  2311 => x"e28d0b80",
  2312 => x"f52d80e2",
  2313 => x"8c0b80f5",
  2314 => x"2d718280",
  2315 => x"290580e2",
  2316 => x"8e0b80f5",
  2317 => x"2d708480",
  2318 => x"80291280",
  2319 => x"e28f0b80",
  2320 => x"f52d7081",
  2321 => x"800a2912",
  2322 => x"7080e894",
  2323 => x"0c80e890",
  2324 => x"08712980",
  2325 => x"e7fc0805",
  2326 => x"7080e880",
  2327 => x"0c80e295",
  2328 => x"0b80f52d",
  2329 => x"80e2940b",
  2330 => x"80f52d71",
  2331 => x"82802905",
  2332 => x"80e2960b",
  2333 => x"80f52d70",
  2334 => x"84808029",
  2335 => x"1280e297",
  2336 => x"0b80f52d",
  2337 => x"70982b81",
  2338 => x"f00a0672",
  2339 => x"057080e8",
  2340 => x"840cfe11",
  2341 => x"7e297705",
  2342 => x"80e8880c",
  2343 => x"52595243",
  2344 => x"545e5152",
  2345 => x"59525d57",
  2346 => x"595780ca",
  2347 => x"860480e1",
  2348 => x"fa0b80f5",
  2349 => x"2d80e1f9",
  2350 => x"0b80f52d",
  2351 => x"71828029",
  2352 => x"057080e7",
  2353 => x"f80c70a0",
  2354 => x"2983ff05",
  2355 => x"70892a70",
  2356 => x"80e88c0c",
  2357 => x"80e1ff0b",
  2358 => x"80f52d80",
  2359 => x"e1fe0b80",
  2360 => x"f52d7182",
  2361 => x"80290570",
  2362 => x"80e8940c",
  2363 => x"7b71291e",
  2364 => x"7080e888",
  2365 => x"0c7d80e8",
  2366 => x"840c7305",
  2367 => x"80e8800c",
  2368 => x"555e5151",
  2369 => x"55558051",
  2370 => x"80c2c92d",
  2371 => x"81557480",
  2372 => x"dfac0c02",
  2373 => x"a8050d04",
  2374 => x"02ec050d",
  2375 => x"7670872c",
  2376 => x"7180ff06",
  2377 => x"55565480",
  2378 => x"e7f4088a",
  2379 => x"3873882c",
  2380 => x"7481ff06",
  2381 => x"545580e1",
  2382 => x"e85280e7",
  2383 => x"fc081551",
  2384 => x"80c0e22d",
  2385 => x"80dfac08",
  2386 => x"5480dfac",
  2387 => x"08802ebb",
  2388 => x"3880e7f4",
  2389 => x"08802e9c",
  2390 => x"38728429",
  2391 => x"80e1e805",
  2392 => x"70085253",
  2393 => x"80d0d22d",
  2394 => x"80dfac08",
  2395 => x"f00a0653",
  2396 => x"80cb8904",
  2397 => x"721080e1",
  2398 => x"e8057080",
  2399 => x"e02d5253",
  2400 => x"80d1832d",
  2401 => x"80dfac08",
  2402 => x"53725473",
  2403 => x"80dfac0c",
  2404 => x"0294050d",
  2405 => x"0402e005",
  2406 => x"0d797084",
  2407 => x"2c80e89c",
  2408 => x"0805718f",
  2409 => x"06525553",
  2410 => x"728b3880",
  2411 => x"e1e85273",
  2412 => x"5180c0e2",
  2413 => x"2d72a029",
  2414 => x"80e1e805",
  2415 => x"54807480",
  2416 => x"f52d5653",
  2417 => x"74732e83",
  2418 => x"38815374",
  2419 => x"81e52e81",
  2420 => x"f5388170",
  2421 => x"74065458",
  2422 => x"72802e81",
  2423 => x"e9388b14",
  2424 => x"80f52d70",
  2425 => x"832a7906",
  2426 => x"5856769c",
  2427 => x"3880ddf0",
  2428 => x"08537289",
  2429 => x"387280e5",
  2430 => x"e80b81b7",
  2431 => x"2d7680dd",
  2432 => x"f00c7353",
  2433 => x"80cdc804",
  2434 => x"758f2e09",
  2435 => x"810681b6",
  2436 => x"38749f06",
  2437 => x"8d2980e5",
  2438 => x"db115153",
  2439 => x"811480f5",
  2440 => x"2d737081",
  2441 => x"055581b7",
  2442 => x"2d831480",
  2443 => x"f52d7370",
  2444 => x"81055581",
  2445 => x"b72d8514",
  2446 => x"80f52d73",
  2447 => x"70810555",
  2448 => x"81b72d87",
  2449 => x"1480f52d",
  2450 => x"73708105",
  2451 => x"5581b72d",
  2452 => x"891480f5",
  2453 => x"2d737081",
  2454 => x"055581b7",
  2455 => x"2d8e1480",
  2456 => x"f52d7370",
  2457 => x"81055581",
  2458 => x"b72d9014",
  2459 => x"80f52d73",
  2460 => x"70810555",
  2461 => x"81b72d92",
  2462 => x"1480f52d",
  2463 => x"73708105",
  2464 => x"5581b72d",
  2465 => x"941480f5",
  2466 => x"2d737081",
  2467 => x"055581b7",
  2468 => x"2d961480",
  2469 => x"f52d7370",
  2470 => x"81055581",
  2471 => x"b72d9814",
  2472 => x"80f52d73",
  2473 => x"70810555",
  2474 => x"81b72d9c",
  2475 => x"1480f52d",
  2476 => x"73708105",
  2477 => x"5581b72d",
  2478 => x"9e1480f5",
  2479 => x"2d7381b7",
  2480 => x"2d7780dd",
  2481 => x"f00c8053",
  2482 => x"7280dfac",
  2483 => x"0c02a005",
  2484 => x"0d0402cc",
  2485 => x"050d7e60",
  2486 => x"5e5a800b",
  2487 => x"80e89808",
  2488 => x"80e89c08",
  2489 => x"595c5680",
  2490 => x"5880e7f8",
  2491 => x"08782e81",
  2492 => x"be38778f",
  2493 => x"06a01757",
  2494 => x"54739238",
  2495 => x"80e1e852",
  2496 => x"76518117",
  2497 => x"5780c0e2",
  2498 => x"2d80e1e8",
  2499 => x"56807680",
  2500 => x"f52d5654",
  2501 => x"74742e83",
  2502 => x"38815474",
  2503 => x"81e52e81",
  2504 => x"82388170",
  2505 => x"7506555c",
  2506 => x"73802e80",
  2507 => x"f6388b16",
  2508 => x"80f52d98",
  2509 => x"06597880",
  2510 => x"ea388b53",
  2511 => x"7c527551",
  2512 => x"80c2882d",
  2513 => x"80dfac08",
  2514 => x"80d9389c",
  2515 => x"16085180",
  2516 => x"d0d22d80",
  2517 => x"dfac0884",
  2518 => x"1b0c9a16",
  2519 => x"80e02d51",
  2520 => x"80d1832d",
  2521 => x"80dfac08",
  2522 => x"80dfac08",
  2523 => x"881c0c80",
  2524 => x"dfac0855",
  2525 => x"5580e7f4",
  2526 => x"08802e9a",
  2527 => x"38941680",
  2528 => x"e02d5180",
  2529 => x"d1832d80",
  2530 => x"dfac0890",
  2531 => x"2b83fff0",
  2532 => x"0a067016",
  2533 => x"51547388",
  2534 => x"1b0c787a",
  2535 => x"0c7b5480",
  2536 => x"cfed0481",
  2537 => x"185880e7",
  2538 => x"f8087826",
  2539 => x"fec43880",
  2540 => x"e7f40880",
  2541 => x"2eb5387a",
  2542 => x"5180ca98",
  2543 => x"2d80dfac",
  2544 => x"0880dfac",
  2545 => x"0880ffff",
  2546 => x"fff80655",
  2547 => x"5b7380ff",
  2548 => x"fffff82e",
  2549 => x"963880df",
  2550 => x"ac08fe05",
  2551 => x"80e7ec08",
  2552 => x"2980e880",
  2553 => x"08055780",
  2554 => x"cde70480",
  2555 => x"547380df",
  2556 => x"ac0c02b4",
  2557 => x"050d0402",
  2558 => x"f4050d74",
  2559 => x"70088105",
  2560 => x"710c7008",
  2561 => x"80e7f008",
  2562 => x"06535371",
  2563 => x"90388813",
  2564 => x"085180ca",
  2565 => x"982d80df",
  2566 => x"ac088814",
  2567 => x"0c810b80",
  2568 => x"dfac0c02",
  2569 => x"8c050d04",
  2570 => x"02f0050d",
  2571 => x"75881108",
  2572 => x"fe0580e7",
  2573 => x"ec082980",
  2574 => x"e8800811",
  2575 => x"720880e7",
  2576 => x"f0080605",
  2577 => x"79555354",
  2578 => x"5480c0e2",
  2579 => x"2d029005",
  2580 => x"0d0402f4",
  2581 => x"050d7470",
  2582 => x"882a83fe",
  2583 => x"80067072",
  2584 => x"982a0772",
  2585 => x"882b87fc",
  2586 => x"80800673",
  2587 => x"982b81f0",
  2588 => x"0a067173",
  2589 => x"070780df",
  2590 => x"ac0c5651",
  2591 => x"5351028c",
  2592 => x"050d0402",
  2593 => x"f8050d02",
  2594 => x"8e0580f5",
  2595 => x"2d74882b",
  2596 => x"077083ff",
  2597 => x"ff0680df",
  2598 => x"ac0c5102",
  2599 => x"88050d04",
  2600 => x"02f4050d",
  2601 => x"74767853",
  2602 => x"54528071",
  2603 => x"25973872",
  2604 => x"70810554",
  2605 => x"80f52d72",
  2606 => x"70810554",
  2607 => x"81b72dff",
  2608 => x"115170eb",
  2609 => x"38807281",
  2610 => x"b72d028c",
  2611 => x"050d0402",
  2612 => x"e8050d77",
  2613 => x"56807056",
  2614 => x"54737624",
  2615 => x"b73880e7",
  2616 => x"f808742e",
  2617 => x"af387351",
  2618 => x"80cb952d",
  2619 => x"80dfac08",
  2620 => x"80dfac08",
  2621 => x"09810570",
  2622 => x"80dfac08",
  2623 => x"079f2a77",
  2624 => x"05811757",
  2625 => x"57535374",
  2626 => x"76248938",
  2627 => x"80e7f808",
  2628 => x"7426d338",
  2629 => x"7280dfac",
  2630 => x"0c029805",
  2631 => x"0d0402f0",
  2632 => x"050d80df",
  2633 => x"a8081651",
  2634 => x"80d1cf2d",
  2635 => x"80dfac08",
  2636 => x"802ea038",
  2637 => x"8b5380df",
  2638 => x"ac085280",
  2639 => x"e5e85180",
  2640 => x"d1a02d80",
  2641 => x"e8a40854",
  2642 => x"73802e87",
  2643 => x"3880e5e8",
  2644 => x"51732d02",
  2645 => x"90050d04",
  2646 => x"02dc050d",
  2647 => x"80705a55",
  2648 => x"7480dfa8",
  2649 => x"0825b538",
  2650 => x"80e7f808",
  2651 => x"752ead38",
  2652 => x"785180cb",
  2653 => x"952d80df",
  2654 => x"ac080981",
  2655 => x"057080df",
  2656 => x"ac08079f",
  2657 => x"2a760581",
  2658 => x"1b5b5654",
  2659 => x"7480dfa8",
  2660 => x"08258938",
  2661 => x"80e7f808",
  2662 => x"7926d538",
  2663 => x"80557880",
  2664 => x"e7f80827",
  2665 => x"81e43878",
  2666 => x"5180cb95",
  2667 => x"2d80dfac",
  2668 => x"08802e81",
  2669 => x"b43880df",
  2670 => x"ac088b05",
  2671 => x"80f52d70",
  2672 => x"842a7081",
  2673 => x"06771078",
  2674 => x"842b80e5",
  2675 => x"e80b80f5",
  2676 => x"2d5c5c53",
  2677 => x"51555673",
  2678 => x"802e80ce",
  2679 => x"38741682",
  2680 => x"2b80d5ae",
  2681 => x"0b80ddfc",
  2682 => x"120c5477",
  2683 => x"75311080",
  2684 => x"e8a81155",
  2685 => x"56907470",
  2686 => x"81055681",
  2687 => x"b72da074",
  2688 => x"81b72d76",
  2689 => x"81ff0681",
  2690 => x"16585473",
  2691 => x"802e8b38",
  2692 => x"9c5380e5",
  2693 => x"e85280d4",
  2694 => x"a1048b53",
  2695 => x"80dfac08",
  2696 => x"5280e8aa",
  2697 => x"165180d4",
  2698 => x"df047416",
  2699 => x"822b80d2",
  2700 => x"9e0b80dd",
  2701 => x"fc120c54",
  2702 => x"7681ff06",
  2703 => x"81165854",
  2704 => x"73802e8b",
  2705 => x"389c5380",
  2706 => x"e5e85280",
  2707 => x"d4d6048b",
  2708 => x"5380dfac",
  2709 => x"08527775",
  2710 => x"311080e8",
  2711 => x"a8055176",
  2712 => x"5580d1a0",
  2713 => x"2d80d4fe",
  2714 => x"04749029",
  2715 => x"75317010",
  2716 => x"80e8a805",
  2717 => x"515480df",
  2718 => x"ac087481",
  2719 => x"b72d8119",
  2720 => x"59748b24",
  2721 => x"a43880d3",
  2722 => x"9e047490",
  2723 => x"29753170",
  2724 => x"1080e8a8",
  2725 => x"058c7731",
  2726 => x"57515480",
  2727 => x"7481b72d",
  2728 => x"9e14ff16",
  2729 => x"565474f3",
  2730 => x"3802a405",
  2731 => x"0d0402fc",
  2732 => x"050d80df",
  2733 => x"a8081351",
  2734 => x"80d1cf2d",
  2735 => x"80dfac08",
  2736 => x"802e8a38",
  2737 => x"80dfac08",
  2738 => x"5180c2c9",
  2739 => x"2d800b80",
  2740 => x"dfa80c80",
  2741 => x"d2d82db0",
  2742 => x"cb2d0284",
  2743 => x"050d0402",
  2744 => x"fc050d72",
  2745 => x"5170fd2e",
  2746 => x"b23870fd",
  2747 => x"248b3870",
  2748 => x"fc2e80d0",
  2749 => x"3880d6ce",
  2750 => x"0470fe2e",
  2751 => x"b93870ff",
  2752 => x"2e098106",
  2753 => x"80c83880",
  2754 => x"dfa80851",
  2755 => x"70802ebe",
  2756 => x"38ff1180",
  2757 => x"dfa80c80",
  2758 => x"d6ce0480",
  2759 => x"dfa808f0",
  2760 => x"057080df",
  2761 => x"a80c5170",
  2762 => x"8025a338",
  2763 => x"800b80df",
  2764 => x"a80c80d6",
  2765 => x"ce0480df",
  2766 => x"a8088105",
  2767 => x"80dfa80c",
  2768 => x"80d6ce04",
  2769 => x"80dfa808",
  2770 => x"900580df",
  2771 => x"a80c80d2",
  2772 => x"d82db0cb",
  2773 => x"2d028405",
  2774 => x"0d0402fc",
  2775 => x"050d800b",
  2776 => x"80dfa80c",
  2777 => x"80d2d82d",
  2778 => x"afc72d80",
  2779 => x"dfac0880",
  2780 => x"df980c80",
  2781 => x"ddf451b1",
  2782 => x"f12d0284",
  2783 => x"050d0471",
  2784 => x"80e8a40c",
  2785 => x"04000000",
  2786 => x"00ffffff",
  2787 => x"ff00ffff",
  2788 => x"ffff00ff",
  2789 => x"ffffff00",
  2790 => x"30313233",
  2791 => x"34353637",
  2792 => x"38394142",
  2793 => x"43444546",
  2794 => x"00000000",
  2795 => x"52657365",
  2796 => x"74000000",
  2797 => x"5363616e",
  2798 => x"6c696e65",
  2799 => x"73000000",
  2800 => x"50414c20",
  2801 => x"2f204e54",
  2802 => x"53430000",
  2803 => x"436f6c6f",
  2804 => x"72000000",
  2805 => x"44696666",
  2806 => x"6963756c",
  2807 => x"74792041",
  2808 => x"00000000",
  2809 => x"44696666",
  2810 => x"6963756c",
  2811 => x"74792042",
  2812 => x"00000000",
  2813 => x"2a537570",
  2814 => x"65726368",
  2815 => x"69702069",
  2816 => x"6e206361",
  2817 => x"72747269",
  2818 => x"64676500",
  2819 => x"2a42616e",
  2820 => x"6b204530",
  2821 => x"00000000",
  2822 => x"2a42616e",
  2823 => x"6b204537",
  2824 => x"00000000",
  2825 => x"53656c65",
  2826 => x"63740000",
  2827 => x"53746172",
  2828 => x"74000000",
  2829 => x"4c6f6164",
  2830 => x"20524f4d",
  2831 => x"20100000",
  2832 => x"45786974",
  2833 => x"00000000",
  2834 => x"524f4d20",
  2835 => x"6c6f6164",
  2836 => x"696e6720",
  2837 => x"6661696c",
  2838 => x"65640000",
  2839 => x"4f4b0000",
  2840 => x"496e6974",
  2841 => x"69616c69",
  2842 => x"7a696e67",
  2843 => x"20534420",
  2844 => x"63617264",
  2845 => x"0a000000",
  2846 => x"436f6c6c",
  2847 => x"6563746f",
  2848 => x"72566973",
  2849 => x"696f6e00",
  2850 => x"64626732",
  2851 => x"00000000",
  2852 => x"16200000",
  2853 => x"14200000",
  2854 => x"15200000",
  2855 => x"53442069",
  2856 => x"6e69742e",
  2857 => x"2e2e0a00",
  2858 => x"53442063",
  2859 => x"61726420",
  2860 => x"72657365",
  2861 => x"74206661",
  2862 => x"696c6564",
  2863 => x"210a0000",
  2864 => x"53444843",
  2865 => x"20657272",
  2866 => x"6f72210a",
  2867 => x"00000000",
  2868 => x"57726974",
  2869 => x"65206661",
  2870 => x"696c6564",
  2871 => x"0a000000",
  2872 => x"52656164",
  2873 => x"20666169",
  2874 => x"6c65640a",
  2875 => x"00000000",
  2876 => x"43617264",
  2877 => x"20696e69",
  2878 => x"74206661",
  2879 => x"696c6564",
  2880 => x"0a000000",
  2881 => x"46415431",
  2882 => x"36202020",
  2883 => x"00000000",
  2884 => x"46415433",
  2885 => x"32202020",
  2886 => x"00000000",
  2887 => x"4e6f2070",
  2888 => x"61727469",
  2889 => x"74696f6e",
  2890 => x"20736967",
  2891 => x"0a000000",
  2892 => x"42616420",
  2893 => x"70617274",
  2894 => x"0a000000",
  2895 => x"4261636b",
  2896 => x"00000000",
  2897 => x"00000002",
  2898 => x"00002b98",
  2899 => x"0000305c",
  2900 => x"00000002",
  2901 => x"00002fd4",
  2902 => x"0000135a",
  2903 => x"00000002",
  2904 => x"00003018",
  2905 => x"00001276",
  2906 => x"00000002",
  2907 => x"00002bac",
  2908 => x"0000035a",
  2909 => x"00000001",
  2910 => x"00002bb4",
  2911 => x"00000000",
  2912 => x"00000001",
  2913 => x"00002bc0",
  2914 => x"00000001",
  2915 => x"00000001",
  2916 => x"00002bcc",
  2917 => x"00000002",
  2918 => x"00000001",
  2919 => x"00002bd4",
  2920 => x"00000003",
  2921 => x"00000001",
  2922 => x"00002be4",
  2923 => x"00000004",
  2924 => x"00000001",
  2925 => x"00002bf4",
  2926 => x"00000005",
  2927 => x"00000001",
  2928 => x"00002c0c",
  2929 => x"00000008",
  2930 => x"00000001",
  2931 => x"00002c18",
  2932 => x"00000009",
  2933 => x"00000002",
  2934 => x"00002c24",
  2935 => x"0000036e",
  2936 => x"00000002",
  2937 => x"00002c2c",
  2938 => x"00000a3f",
  2939 => x"00000002",
  2940 => x"00002c34",
  2941 => x"00002b5a",
  2942 => x"00000002",
  2943 => x"00002c40",
  2944 => x"000017e4",
  2945 => x"00000000",
  2946 => x"00000000",
  2947 => x"00000000",
  2948 => x"00000004",
  2949 => x"00002c48",
  2950 => x"00002e10",
  2951 => x"00000004",
  2952 => x"00002c5c",
  2953 => x"00002d50",
  2954 => x"00000000",
  2955 => x"00000000",
  2956 => x"00000000",
  2957 => x"00000000",
  2958 => x"00000000",
  2959 => x"00000000",
  2960 => x"00000000",
  2961 => x"00000000",
  2962 => x"00000000",
  2963 => x"00000000",
  2964 => x"00000000",
  2965 => x"00000000",
  2966 => x"00000000",
  2967 => x"00000000",
  2968 => x"00000000",
  2969 => x"00000000",
  2970 => x"00000000",
  2971 => x"00000000",
  2972 => x"00000000",
  2973 => x"00000000",
  2974 => x"76f55a1c",
  2975 => x"f21c051c",
  2976 => x"1c1c1c1c",
  2977 => x"f2f5ebf4",
  2978 => x"5a000000",
  2979 => x"00000000",
  2980 => x"00000000",
  2981 => x"00000000",
  2982 => x"00000000",
  2983 => x"00000000",
  2984 => x"00000000",
  2985 => x"00000000",
  2986 => x"00000000",
  2987 => x"00000000",
  2988 => x"00000000",
  2989 => x"00000000",
  2990 => x"00000000",
  2991 => x"00000000",
  2992 => x"00000000",
  2993 => x"00000000",
  2994 => x"00000000",
  2995 => x"00000000",
  2996 => x"00000000",
  2997 => x"0001ffff",
  2998 => x"0001ffff",
  2999 => x"0001ffff",
  3000 => x"00000000",
  3001 => x"00000000",
  3002 => x"00000006",
  3003 => x"00000000",
  3004 => x"00000000",
  3005 => x"00000002",
  3006 => x"00003428",
  3007 => x"0000291e",
  3008 => x"00000002",
  3009 => x"00003446",
  3010 => x"0000291e",
  3011 => x"00000002",
  3012 => x"00003464",
  3013 => x"0000291e",
  3014 => x"00000002",
  3015 => x"00003482",
  3016 => x"0000291e",
  3017 => x"00000002",
  3018 => x"000034a0",
  3019 => x"0000291e",
  3020 => x"00000002",
  3021 => x"000034be",
  3022 => x"0000291e",
  3023 => x"00000002",
  3024 => x"000034dc",
  3025 => x"0000291e",
  3026 => x"00000002",
  3027 => x"000034fa",
  3028 => x"0000291e",
  3029 => x"00000002",
  3030 => x"00003518",
  3031 => x"0000291e",
  3032 => x"00000002",
  3033 => x"00003536",
  3034 => x"0000291e",
  3035 => x"00000002",
  3036 => x"00003554",
  3037 => x"0000291e",
  3038 => x"00000002",
  3039 => x"00003572",
  3040 => x"0000291e",
  3041 => x"00000002",
  3042 => x"00003590",
  3043 => x"0000291e",
  3044 => x"00000004",
  3045 => x"00002d3c",
  3046 => x"00000000",
  3047 => x"00000000",
  3048 => x"00000000",
  3049 => x"00002adf",
  3050 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

