-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80e1",
     9 => x"b8080b0b",
    10 => x"80e1bc08",
    11 => x"0b0b80e1",
    12 => x"c0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"e1c00c0b",
    16 => x"0b80e1bc",
    17 => x"0c0b0b80",
    18 => x"e1b80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d8f0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80e1b870",
    57 => x"80ecf027",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a6d9",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80e1",
    65 => x"c80c9f0b",
    66 => x"80e1cc0c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"e1cc08ff",
    70 => x"0580e1cc",
    71 => x"0c80e1cc",
    72 => x"088025e8",
    73 => x"3880e1c8",
    74 => x"08ff0580",
    75 => x"e1c80c80",
    76 => x"e1c80880",
    77 => x"25d03880",
    78 => x"0b80e1cc",
    79 => x"0c800b80",
    80 => x"e1c80c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80e1c808",
   100 => x"25913882",
   101 => x"c82d80e1",
   102 => x"c808ff05",
   103 => x"80e1c80c",
   104 => x"838a0480",
   105 => x"e1c80880",
   106 => x"e1cc0853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80e1c808",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"e1cc0881",
   116 => x"0580e1cc",
   117 => x"0c80e1cc",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80e1cc",
   121 => x"0c80e1c8",
   122 => x"08810580",
   123 => x"e1c80c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480e1",
   128 => x"cc088105",
   129 => x"80e1cc0c",
   130 => x"80e1cc08",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80e1cc",
   134 => x"0c80e1c8",
   135 => x"08810580",
   136 => x"e1c80c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"e1d00cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"e1d00c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280e1",
   177 => x"d0088407",
   178 => x"80e1d00c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80dc",
   183 => x"c40c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80e1d0",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80e1",
   208 => x"b80c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02f4050d",
  1093 => x"74765452",
  1094 => x"72708105",
  1095 => x"5480f52d",
  1096 => x"51707270",
  1097 => x"81055481",
  1098 => x"b72d70ec",
  1099 => x"38707281",
  1100 => x"b72d028c",
  1101 => x"050d0402",
  1102 => x"f4050d80",
  1103 => x"dce00b80",
  1104 => x"f52d80df",
  1105 => x"c8087081",
  1106 => x"06535452",
  1107 => x"70802e85",
  1108 => x"38718407",
  1109 => x"5272812a",
  1110 => x"70810651",
  1111 => x"5170802e",
  1112 => x"85387182",
  1113 => x"07527282",
  1114 => x"2a708106",
  1115 => x"51517080",
  1116 => x"2e853871",
  1117 => x"81075272",
  1118 => x"832a7081",
  1119 => x"06515170",
  1120 => x"802e8538",
  1121 => x"71880752",
  1122 => x"72842a70",
  1123 => x"81065151",
  1124 => x"70802e85",
  1125 => x"38719007",
  1126 => x"5272852a",
  1127 => x"70810651",
  1128 => x"5170802e",
  1129 => x"853871a0",
  1130 => x"07527288",
  1131 => x"2a708106",
  1132 => x"51517080",
  1133 => x"2e863871",
  1134 => x"80c00752",
  1135 => x"72892a70",
  1136 => x"81065151",
  1137 => x"70802e86",
  1138 => x"38718180",
  1139 => x"075271fc",
  1140 => x"0c7180e1",
  1141 => x"b80c028c",
  1142 => x"050d0402",
  1143 => x"cc050d7e",
  1144 => x"5d800b80",
  1145 => x"dfc80881",
  1146 => x"8006715c",
  1147 => x"5d5b810b",
  1148 => x"ec0c840b",
  1149 => x"ec0c7c52",
  1150 => x"80e1d451",
  1151 => x"80ce932d",
  1152 => x"80e1b808",
  1153 => x"7b2e80ff",
  1154 => x"3880e1d8",
  1155 => x"087bff12",
  1156 => x"57595774",
  1157 => x"7b2e8b38",
  1158 => x"81187581",
  1159 => x"2a565874",
  1160 => x"f738f718",
  1161 => x"58815b80",
  1162 => x"772580db",
  1163 => x"38775274",
  1164 => x"5184a82d",
  1165 => x"80e2a852",
  1166 => x"80e1d451",
  1167 => x"80d0e82d",
  1168 => x"80e1b808",
  1169 => x"802ea638",
  1170 => x"80e2a859",
  1171 => x"7ba73883",
  1172 => x"ff567870",
  1173 => x"81055a80",
  1174 => x"f52d7a81",
  1175 => x"1c5ce40c",
  1176 => x"e80cff16",
  1177 => x"56758025",
  1178 => x"e938a4f5",
  1179 => x"0480e1b8",
  1180 => x"085b8480",
  1181 => x"5780e1d4",
  1182 => x"5180d0b7",
  1183 => x"2dfc8017",
  1184 => x"81165657",
  1185 => x"a4a70480",
  1186 => x"e1d808f8",
  1187 => x"0c881d54",
  1188 => x"807480f5",
  1189 => x"2d7081ff",
  1190 => x"06555855",
  1191 => x"72752eb6",
  1192 => x"38811480",
  1193 => x"f52d5372",
  1194 => x"752eab38",
  1195 => x"74821580",
  1196 => x"f52d5456",
  1197 => x"7280d32e",
  1198 => x"09810683",
  1199 => x"38815672",
  1200 => x"80f33270",
  1201 => x"09810570",
  1202 => x"80257807",
  1203 => x"51515372",
  1204 => x"802e8338",
  1205 => x"a0558077",
  1206 => x"81ff0654",
  1207 => x"567280c5",
  1208 => x"2e098106",
  1209 => x"83388156",
  1210 => x"7280e532",
  1211 => x"70098105",
  1212 => x"70802578",
  1213 => x"07515153",
  1214 => x"72802ea4",
  1215 => x"38811480",
  1216 => x"f52d5372",
  1217 => x"b02e0981",
  1218 => x"06893874",
  1219 => x"82800755",
  1220 => x"a6a00472",
  1221 => x"b72e0981",
  1222 => x"06863874",
  1223 => x"84800755",
  1224 => x"80dfc808",
  1225 => x"f9df0675",
  1226 => x"0780dfc8",
  1227 => x"0ca2b72d",
  1228 => x"800be00c",
  1229 => x"805186da",
  1230 => x"2d86c72d",
  1231 => x"7a802e88",
  1232 => x"3880dccc",
  1233 => x"51a6cc04",
  1234 => x"80ddf451",
  1235 => x"b0dc2d7a",
  1236 => x"80e1b80c",
  1237 => x"02b4050d",
  1238 => x"0402f405",
  1239 => x"0d840bec",
  1240 => x"0c810be0",
  1241 => x"0cae992d",
  1242 => x"a7f32d81",
  1243 => x"f92d8352",
  1244 => x"adfc2d81",
  1245 => x"51858d2d",
  1246 => x"ff125271",
  1247 => x"8025f138",
  1248 => x"840bec0c",
  1249 => x"80dac851",
  1250 => x"86a02d80",
  1251 => x"c2ef2d80",
  1252 => x"e1b80880",
  1253 => x"2e80c538",
  1254 => x"80dae051",
  1255 => x"86a02da3",
  1256 => x"db5180d8",
  1257 => x"e82d80dc",
  1258 => x"cc51b0dc",
  1259 => x"2daebb2d",
  1260 => x"a99e2d80",
  1261 => x"e1b80881",
  1262 => x"06527180",
  1263 => x"2e863880",
  1264 => x"5194bf2d",
  1265 => x"b0ef2d80",
  1266 => x"e1b80852",
  1267 => x"a2b72d86",
  1268 => x"53718338",
  1269 => x"845372ec",
  1270 => x"0ca7b004",
  1271 => x"800b80e1",
  1272 => x"b80c028c",
  1273 => x"050d0471",
  1274 => x"980c04ff",
  1275 => x"b00880e1",
  1276 => x"b80c0481",
  1277 => x"0bffb00c",
  1278 => x"04800bff",
  1279 => x"b00c0402",
  1280 => x"d8050dff",
  1281 => x"b40887ff",
  1282 => x"ff065a81",
  1283 => x"54807080",
  1284 => x"dfb40880",
  1285 => x"dfb80880",
  1286 => x"df905b59",
  1287 => x"575a5879",
  1288 => x"74067575",
  1289 => x"06525271",
  1290 => x"712e8d38",
  1291 => x"8077818a",
  1292 => x"2d730975",
  1293 => x"06720755",
  1294 => x"7680e02d",
  1295 => x"7083ffff",
  1296 => x"06535171",
  1297 => x"80e42e09",
  1298 => x"8106a238",
  1299 => x"74740670",
  1300 => x"77760632",
  1301 => x"70098105",
  1302 => x"7072079f",
  1303 => x"2a7b0577",
  1304 => x"097a0674",
  1305 => x"075a5b53",
  1306 => x"5353a8fb",
  1307 => x"047180e4",
  1308 => x"26893881",
  1309 => x"11517077",
  1310 => x"818a2d73",
  1311 => x"10811a82",
  1312 => x"19595a54",
  1313 => x"907925ff",
  1314 => x"96387580",
  1315 => x"dfb80c74",
  1316 => x"80dfb40c",
  1317 => x"7780e1b8",
  1318 => x"0c02a805",
  1319 => x"0d0402d0",
  1320 => x"050d805c",
  1321 => x"aaae0480",
  1322 => x"e1b80881",
  1323 => x"f02e0981",
  1324 => x"068a3881",
  1325 => x"0b80dfc0",
  1326 => x"0caaae04",
  1327 => x"80e1b808",
  1328 => x"81e02e09",
  1329 => x"81068a38",
  1330 => x"810b80df",
  1331 => x"c40caaae",
  1332 => x"0480e1b8",
  1333 => x"085280df",
  1334 => x"c408802e",
  1335 => x"893880e1",
  1336 => x"b8088180",
  1337 => x"05527184",
  1338 => x"2c728f06",
  1339 => x"535380df",
  1340 => x"c008802e",
  1341 => x"9a387284",
  1342 => x"2980de98",
  1343 => x"05721381",
  1344 => x"712b7009",
  1345 => x"73080673",
  1346 => x"0c515353",
  1347 => x"aaa20472",
  1348 => x"842980de",
  1349 => x"98057213",
  1350 => x"83712b72",
  1351 => x"0807720c",
  1352 => x"5353800b",
  1353 => x"80dfc40c",
  1354 => x"800b80df",
  1355 => x"c00c80e1",
  1356 => x"e051acef",
  1357 => x"2d80e1b8",
  1358 => x"08ff24fe",
  1359 => x"ea38a7ff",
  1360 => x"2d80e1b8",
  1361 => x"08802e81",
  1362 => x"b0388159",
  1363 => x"800b80df",
  1364 => x"bc0880df",
  1365 => x"b80880de",
  1366 => x"ec5a5c5c",
  1367 => x"587a7906",
  1368 => x"7a7a0654",
  1369 => x"5271732e",
  1370 => x"80f83872",
  1371 => x"09810570",
  1372 => x"74078025",
  1373 => x"80ded81a",
  1374 => x"80f52d70",
  1375 => x"842c718f",
  1376 => x"06585357",
  1377 => x"57527580",
  1378 => x"2ea33871",
  1379 => x"842980de",
  1380 => x"98057415",
  1381 => x"83712b72",
  1382 => x"0807720c",
  1383 => x"54527680",
  1384 => x"e02d8105",
  1385 => x"52717781",
  1386 => x"8a2dabc3",
  1387 => x"04718429",
  1388 => x"80de9805",
  1389 => x"74158171",
  1390 => x"2b700973",
  1391 => x"0806730c",
  1392 => x"51535374",
  1393 => x"85327009",
  1394 => x"81057080",
  1395 => x"25515152",
  1396 => x"75802e8e",
  1397 => x"38817073",
  1398 => x"06535371",
  1399 => x"802e8338",
  1400 => x"725c7810",
  1401 => x"81198219",
  1402 => x"59595990",
  1403 => x"7825feed",
  1404 => x"3880dfb8",
  1405 => x"0880dfbc",
  1406 => x"0c7b80e1",
  1407 => x"b80c02b0",
  1408 => x"050d0402",
  1409 => x"f8050d80",
  1410 => x"de98528f",
  1411 => x"51807270",
  1412 => x"8405540c",
  1413 => x"ff115170",
  1414 => x"8025f238",
  1415 => x"0288050d",
  1416 => x"0402f005",
  1417 => x"0d7551a7",
  1418 => x"f92d7082",
  1419 => x"2cfc0680",
  1420 => x"de981172",
  1421 => x"109e0671",
  1422 => x"0870722a",
  1423 => x"70830682",
  1424 => x"742b7009",
  1425 => x"7406760c",
  1426 => x"54515657",
  1427 => x"535153a7",
  1428 => x"f32d7180",
  1429 => x"e1b80c02",
  1430 => x"90050d04",
  1431 => x"02fc050d",
  1432 => x"72518071",
  1433 => x"0c800b84",
  1434 => x"120c0284",
  1435 => x"050d0402",
  1436 => x"f0050d75",
  1437 => x"70088412",
  1438 => x"08535353",
  1439 => x"ff547171",
  1440 => x"2ea838a7",
  1441 => x"f92d8413",
  1442 => x"08708429",
  1443 => x"14881170",
  1444 => x"087081ff",
  1445 => x"06841808",
  1446 => x"81118706",
  1447 => x"841a0c53",
  1448 => x"51555151",
  1449 => x"51a7f32d",
  1450 => x"71547380",
  1451 => x"e1b80c02",
  1452 => x"90050d04",
  1453 => x"02f8050d",
  1454 => x"a7f92de0",
  1455 => x"08708b2a",
  1456 => x"70810651",
  1457 => x"52527080",
  1458 => x"2ea13880",
  1459 => x"e1e00870",
  1460 => x"842980e1",
  1461 => x"e8057381",
  1462 => x"ff06710c",
  1463 => x"515180e1",
  1464 => x"e0088111",
  1465 => x"870680e1",
  1466 => x"e00c5180",
  1467 => x"0b80e288",
  1468 => x"0ca7eb2d",
  1469 => x"a7f32d02",
  1470 => x"88050d04",
  1471 => x"02fc050d",
  1472 => x"a7f92d81",
  1473 => x"0b80e288",
  1474 => x"0ca7f32d",
  1475 => x"80e28808",
  1476 => x"5170f938",
  1477 => x"0284050d",
  1478 => x"0402fc05",
  1479 => x"0d80e1e0",
  1480 => x"51acdc2d",
  1481 => x"ac832dad",
  1482 => x"b451a7e7",
  1483 => x"2d028405",
  1484 => x"0d0480e2",
  1485 => x"940880e1",
  1486 => x"b80c0402",
  1487 => x"fc050d81",
  1488 => x"0b80dfcc",
  1489 => x"0c815185",
  1490 => x"8d2d0284",
  1491 => x"050d0402",
  1492 => x"fc050dae",
  1493 => x"d904a99e",
  1494 => x"2d80f651",
  1495 => x"aca12d80",
  1496 => x"e1b808f2",
  1497 => x"3880da51",
  1498 => x"aca12d80",
  1499 => x"e1b808e6",
  1500 => x"3880e1b8",
  1501 => x"0880dfcc",
  1502 => x"0c80e1b8",
  1503 => x"0851858d",
  1504 => x"2d028405",
  1505 => x"0d0402ec",
  1506 => x"050d7654",
  1507 => x"8052870b",
  1508 => x"881580f5",
  1509 => x"2d565374",
  1510 => x"72248338",
  1511 => x"a0537251",
  1512 => x"83842d81",
  1513 => x"128b1580",
  1514 => x"f52d5452",
  1515 => x"727225de",
  1516 => x"38029405",
  1517 => x"0d0402f0",
  1518 => x"050d80e2",
  1519 => x"94085481",
  1520 => x"f92d800b",
  1521 => x"80e2980c",
  1522 => x"7308802e",
  1523 => x"81893882",
  1524 => x"0b80e1cc",
  1525 => x"0c80e298",
  1526 => x"088f0680",
  1527 => x"e1c80c73",
  1528 => x"08527183",
  1529 => x"2e963871",
  1530 => x"83268938",
  1531 => x"71812eb0",
  1532 => x"38b0c004",
  1533 => x"71852ea0",
  1534 => x"38b0c004",
  1535 => x"881480f5",
  1536 => x"2d841508",
  1537 => x"80daf853",
  1538 => x"545286a0",
  1539 => x"2d718429",
  1540 => x"13700852",
  1541 => x"52b0c404",
  1542 => x"7351af86",
  1543 => x"2db0c004",
  1544 => x"80dfc808",
  1545 => x"8815082c",
  1546 => x"70810651",
  1547 => x"5271802e",
  1548 => x"883880da",
  1549 => x"fc51b0bd",
  1550 => x"0480db80",
  1551 => x"5186a02d",
  1552 => x"84140851",
  1553 => x"86a02d80",
  1554 => x"e2980881",
  1555 => x"0580e298",
  1556 => x"0c8c1454",
  1557 => x"afc80402",
  1558 => x"90050d04",
  1559 => x"7180e294",
  1560 => x"0cafb62d",
  1561 => x"80e29808",
  1562 => x"ff0580e2",
  1563 => x"9c0c0402",
  1564 => x"e8050d80",
  1565 => x"e2940880",
  1566 => x"e2a00857",
  1567 => x"5580f651",
  1568 => x"aca12d80",
  1569 => x"e1b80881",
  1570 => x"2a708106",
  1571 => x"51527180",
  1572 => x"2ea438b1",
  1573 => x"9904a99e",
  1574 => x"2d80f651",
  1575 => x"aca12d80",
  1576 => x"e1b808f2",
  1577 => x"3880dfcc",
  1578 => x"08813270",
  1579 => x"80dfcc0c",
  1580 => x"70525285",
  1581 => x"8d2d800b",
  1582 => x"80e28c0c",
  1583 => x"800b80e2",
  1584 => x"900c80df",
  1585 => x"cc08838d",
  1586 => x"3880da51",
  1587 => x"aca12d80",
  1588 => x"e1b80880",
  1589 => x"2e8c3880",
  1590 => x"e28c0881",
  1591 => x"800780e2",
  1592 => x"8c0c80d9",
  1593 => x"51aca12d",
  1594 => x"80e1b808",
  1595 => x"802e8c38",
  1596 => x"80e28c08",
  1597 => x"80c00780",
  1598 => x"e28c0c81",
  1599 => x"9451aca1",
  1600 => x"2d80e1b8",
  1601 => x"08802e8b",
  1602 => x"3880e28c",
  1603 => x"08900780",
  1604 => x"e28c0c81",
  1605 => x"9151aca1",
  1606 => x"2d80e1b8",
  1607 => x"08802e8b",
  1608 => x"3880e28c",
  1609 => x"08a00780",
  1610 => x"e28c0c81",
  1611 => x"f551aca1",
  1612 => x"2d80e1b8",
  1613 => x"08802e8b",
  1614 => x"3880e28c",
  1615 => x"08810780",
  1616 => x"e28c0c81",
  1617 => x"f251aca1",
  1618 => x"2d80e1b8",
  1619 => x"08802e8b",
  1620 => x"3880e28c",
  1621 => x"08820780",
  1622 => x"e28c0c81",
  1623 => x"eb51aca1",
  1624 => x"2d80e1b8",
  1625 => x"08802e8b",
  1626 => x"3880e28c",
  1627 => x"08840780",
  1628 => x"e28c0c81",
  1629 => x"f451aca1",
  1630 => x"2d80e1b8",
  1631 => x"08802e8b",
  1632 => x"3880e28c",
  1633 => x"08880780",
  1634 => x"e28c0c80",
  1635 => x"d851aca1",
  1636 => x"2d80e1b8",
  1637 => x"08802e8c",
  1638 => x"3880e290",
  1639 => x"08818007",
  1640 => x"80e2900c",
  1641 => x"9251aca1",
  1642 => x"2d80e1b8",
  1643 => x"08802e8c",
  1644 => x"3880e290",
  1645 => x"0880c007",
  1646 => x"80e2900c",
  1647 => x"9451aca1",
  1648 => x"2d80e1b8",
  1649 => x"08802e8b",
  1650 => x"3880e290",
  1651 => x"08900780",
  1652 => x"e2900c91",
  1653 => x"51aca12d",
  1654 => x"80e1b808",
  1655 => x"802e8b38",
  1656 => x"80e29008",
  1657 => x"a00780e2",
  1658 => x"900c9d51",
  1659 => x"aca12d80",
  1660 => x"e1b80880",
  1661 => x"2e8b3880",
  1662 => x"e2900881",
  1663 => x"0780e290",
  1664 => x"0c9b51ac",
  1665 => x"a12d80e1",
  1666 => x"b808802e",
  1667 => x"8b3880e2",
  1668 => x"90088207",
  1669 => x"80e2900c",
  1670 => x"9c51aca1",
  1671 => x"2d80e1b8",
  1672 => x"08802e8b",
  1673 => x"3880e290",
  1674 => x"08840780",
  1675 => x"e2900ca3",
  1676 => x"51aca12d",
  1677 => x"80e1b808",
  1678 => x"802e8b38",
  1679 => x"80e29008",
  1680 => x"880780e2",
  1681 => x"900c81fd",
  1682 => x"51aca12d",
  1683 => x"81fa51ac",
  1684 => x"a12dbaaa",
  1685 => x"0481f551",
  1686 => x"aca12d80",
  1687 => x"e1b80881",
  1688 => x"2a708106",
  1689 => x"51527180",
  1690 => x"2eb33880",
  1691 => x"e29c0852",
  1692 => x"71802e8a",
  1693 => x"38ff1280",
  1694 => x"e29c0cb5",
  1695 => x"9d0480e2",
  1696 => x"98081080",
  1697 => x"e2980805",
  1698 => x"70842916",
  1699 => x"51528812",
  1700 => x"08802e89",
  1701 => x"38ff5188",
  1702 => x"12085271",
  1703 => x"2d81f251",
  1704 => x"aca12d80",
  1705 => x"e1b80881",
  1706 => x"2a708106",
  1707 => x"51527180",
  1708 => x"2eb43880",
  1709 => x"e29808ff",
  1710 => x"1180e29c",
  1711 => x"08565353",
  1712 => x"7372258a",
  1713 => x"38811480",
  1714 => x"e29c0cb5",
  1715 => x"e6047210",
  1716 => x"13708429",
  1717 => x"16515288",
  1718 => x"1208802e",
  1719 => x"8938fe51",
  1720 => x"88120852",
  1721 => x"712d81fd",
  1722 => x"51aca12d",
  1723 => x"80e1b808",
  1724 => x"812a7081",
  1725 => x"06515271",
  1726 => x"802eb138",
  1727 => x"80e29c08",
  1728 => x"802e8a38",
  1729 => x"800b80e2",
  1730 => x"9c0cb6ac",
  1731 => x"0480e298",
  1732 => x"081080e2",
  1733 => x"98080570",
  1734 => x"84291651",
  1735 => x"52881208",
  1736 => x"802e8938",
  1737 => x"fd518812",
  1738 => x"0852712d",
  1739 => x"81fa51ac",
  1740 => x"a12d80e1",
  1741 => x"b808812a",
  1742 => x"70810651",
  1743 => x"5271802e",
  1744 => x"b13880e2",
  1745 => x"9808ff11",
  1746 => x"545280e2",
  1747 => x"9c087325",
  1748 => x"89387280",
  1749 => x"e29c0cb6",
  1750 => x"f2047110",
  1751 => x"12708429",
  1752 => x"16515288",
  1753 => x"1208802e",
  1754 => x"8938fc51",
  1755 => x"88120852",
  1756 => x"712d80e2",
  1757 => x"9c087053",
  1758 => x"5473802e",
  1759 => x"8a388c15",
  1760 => x"ff155555",
  1761 => x"b6f90482",
  1762 => x"0b80e1cc",
  1763 => x"0c718f06",
  1764 => x"80e1c80c",
  1765 => x"81eb51ac",
  1766 => x"a12d80e1",
  1767 => x"b808812a",
  1768 => x"70810651",
  1769 => x"5271802e",
  1770 => x"ad387408",
  1771 => x"852e0981",
  1772 => x"06a43888",
  1773 => x"1580f52d",
  1774 => x"ff055271",
  1775 => x"881681b7",
  1776 => x"2d71982b",
  1777 => x"52718025",
  1778 => x"8838800b",
  1779 => x"881681b7",
  1780 => x"2d7451af",
  1781 => x"862d81f4",
  1782 => x"51aca12d",
  1783 => x"80e1b808",
  1784 => x"812a7081",
  1785 => x"06515271",
  1786 => x"802eb338",
  1787 => x"7408852e",
  1788 => x"098106aa",
  1789 => x"38881580",
  1790 => x"f52d8105",
  1791 => x"52718816",
  1792 => x"81b72d71",
  1793 => x"81ff068b",
  1794 => x"1680f52d",
  1795 => x"54527272",
  1796 => x"27873872",
  1797 => x"881681b7",
  1798 => x"2d7451af",
  1799 => x"862d80da",
  1800 => x"51aca12d",
  1801 => x"80e1b808",
  1802 => x"812a7081",
  1803 => x"06515271",
  1804 => x"802e81ad",
  1805 => x"3880e294",
  1806 => x"0880e29c",
  1807 => x"08555373",
  1808 => x"802e8a38",
  1809 => x"8c13ff15",
  1810 => x"5553b8bf",
  1811 => x"04720852",
  1812 => x"71822ea6",
  1813 => x"38718226",
  1814 => x"89387181",
  1815 => x"2eaa38b9",
  1816 => x"e1047183",
  1817 => x"2eb43871",
  1818 => x"842e0981",
  1819 => x"0680f238",
  1820 => x"88130851",
  1821 => x"b0dc2db9",
  1822 => x"e10480e2",
  1823 => x"9c085188",
  1824 => x"13085271",
  1825 => x"2db9e104",
  1826 => x"810b8814",
  1827 => x"082b80df",
  1828 => x"c8083280",
  1829 => x"dfc80cb9",
  1830 => x"b5048813",
  1831 => x"80f52d81",
  1832 => x"058b1480",
  1833 => x"f52d5354",
  1834 => x"71742483",
  1835 => x"38805473",
  1836 => x"881481b7",
  1837 => x"2dafb62d",
  1838 => x"b9e10475",
  1839 => x"08802ea4",
  1840 => x"38750851",
  1841 => x"aca12d80",
  1842 => x"e1b80881",
  1843 => x"06527180",
  1844 => x"2e8c3880",
  1845 => x"e29c0851",
  1846 => x"84160852",
  1847 => x"712d8816",
  1848 => x"5675d838",
  1849 => x"8054800b",
  1850 => x"80e1cc0c",
  1851 => x"738f0680",
  1852 => x"e1c80ca0",
  1853 => x"527380e2",
  1854 => x"9c082e09",
  1855 => x"81069938",
  1856 => x"80e29808",
  1857 => x"ff057432",
  1858 => x"70098105",
  1859 => x"7072079f",
  1860 => x"2a917131",
  1861 => x"51515353",
  1862 => x"71518384",
  1863 => x"2d811454",
  1864 => x"8e7425c2",
  1865 => x"3880dfcc",
  1866 => x"08527180",
  1867 => x"e1b80c02",
  1868 => x"98050d04",
  1869 => x"02f4050d",
  1870 => x"d45281ff",
  1871 => x"720c7108",
  1872 => x"5381ff72",
  1873 => x"0c72882b",
  1874 => x"83fe8006",
  1875 => x"72087081",
  1876 => x"ff065152",
  1877 => x"5381ff72",
  1878 => x"0c727107",
  1879 => x"882b7208",
  1880 => x"7081ff06",
  1881 => x"51525381",
  1882 => x"ff720c72",
  1883 => x"7107882b",
  1884 => x"72087081",
  1885 => x"ff067207",
  1886 => x"80e1b80c",
  1887 => x"5253028c",
  1888 => x"050d0402",
  1889 => x"f4050d74",
  1890 => x"767181ff",
  1891 => x"06d40c53",
  1892 => x"5380e2a4",
  1893 => x"08853871",
  1894 => x"892b5271",
  1895 => x"982ad40c",
  1896 => x"71902a70",
  1897 => x"81ff06d4",
  1898 => x"0c517188",
  1899 => x"2a7081ff",
  1900 => x"06d40c51",
  1901 => x"7181ff06",
  1902 => x"d40c7290",
  1903 => x"2a7081ff",
  1904 => x"06d40c51",
  1905 => x"d4087081",
  1906 => x"ff065151",
  1907 => x"82b8bf52",
  1908 => x"7081ff2e",
  1909 => x"09810694",
  1910 => x"3881ff0b",
  1911 => x"d40cd408",
  1912 => x"7081ff06",
  1913 => x"ff145451",
  1914 => x"5171e538",
  1915 => x"7080e1b8",
  1916 => x"0c028c05",
  1917 => x"0d0402fc",
  1918 => x"050d81c7",
  1919 => x"5181ff0b",
  1920 => x"d40cff11",
  1921 => x"51708025",
  1922 => x"f4380284",
  1923 => x"050d0402",
  1924 => x"f4050d81",
  1925 => x"ff0bd40c",
  1926 => x"93538052",
  1927 => x"87fc80c1",
  1928 => x"51bb832d",
  1929 => x"80e1b808",
  1930 => x"8b3881ff",
  1931 => x"0bd40c81",
  1932 => x"53bcbd04",
  1933 => x"bbf62dff",
  1934 => x"135372de",
  1935 => x"387280e1",
  1936 => x"b80c028c",
  1937 => x"050d0402",
  1938 => x"ec050d81",
  1939 => x"0b80e2a4",
  1940 => x"0c8454d0",
  1941 => x"08708f2a",
  1942 => x"70810651",
  1943 => x"515372f3",
  1944 => x"3872d00c",
  1945 => x"bbf62d80",
  1946 => x"db845186",
  1947 => x"a02dd008",
  1948 => x"708f2a70",
  1949 => x"81065151",
  1950 => x"5372f338",
  1951 => x"810bd00c",
  1952 => x"b1538052",
  1953 => x"84d480c0",
  1954 => x"51bb832d",
  1955 => x"80e1b808",
  1956 => x"812e9338",
  1957 => x"72822ebf",
  1958 => x"38ff1353",
  1959 => x"72e438ff",
  1960 => x"145473ff",
  1961 => x"ae38bbf6",
  1962 => x"2d83aa52",
  1963 => x"849c80c8",
  1964 => x"51bb832d",
  1965 => x"80e1b808",
  1966 => x"812e0981",
  1967 => x"069338ba",
  1968 => x"b42d80e1",
  1969 => x"b80883ff",
  1970 => x"ff065372",
  1971 => x"83aa2e9f",
  1972 => x"38bc8f2d",
  1973 => x"bdea0480",
  1974 => x"db905186",
  1975 => x"a02d8053",
  1976 => x"bfbf0480",
  1977 => x"dba85186",
  1978 => x"a02d8054",
  1979 => x"bf900481",
  1980 => x"ff0bd40c",
  1981 => x"b154bbf6",
  1982 => x"2d8fcf53",
  1983 => x"805287fc",
  1984 => x"80f751bb",
  1985 => x"832d80e1",
  1986 => x"b8085580",
  1987 => x"e1b80881",
  1988 => x"2e098106",
  1989 => x"9c3881ff",
  1990 => x"0bd40c82",
  1991 => x"0a52849c",
  1992 => x"80e951bb",
  1993 => x"832d80e1",
  1994 => x"b808802e",
  1995 => x"8d38bbf6",
  1996 => x"2dff1353",
  1997 => x"72c638bf",
  1998 => x"830481ff",
  1999 => x"0bd40c80",
  2000 => x"e1b80852",
  2001 => x"87fc80fa",
  2002 => x"51bb832d",
  2003 => x"80e1b808",
  2004 => x"b23881ff",
  2005 => x"0bd40cd4",
  2006 => x"085381ff",
  2007 => x"0bd40c81",
  2008 => x"ff0bd40c",
  2009 => x"81ff0bd4",
  2010 => x"0c81ff0b",
  2011 => x"d40c7286",
  2012 => x"2a708106",
  2013 => x"76565153",
  2014 => x"72963880",
  2015 => x"e1b80854",
  2016 => x"bf900473",
  2017 => x"822efedb",
  2018 => x"38ff1454",
  2019 => x"73fee738",
  2020 => x"7380e2a4",
  2021 => x"0c738b38",
  2022 => x"815287fc",
  2023 => x"80d051bb",
  2024 => x"832d81ff",
  2025 => x"0bd40cd0",
  2026 => x"08708f2a",
  2027 => x"70810651",
  2028 => x"515372f3",
  2029 => x"3872d00c",
  2030 => x"81ff0bd4",
  2031 => x"0c815372",
  2032 => x"80e1b80c",
  2033 => x"0294050d",
  2034 => x"0402e805",
  2035 => x"0d785580",
  2036 => x"5681ff0b",
  2037 => x"d40cd008",
  2038 => x"708f2a70",
  2039 => x"81065151",
  2040 => x"5372f338",
  2041 => x"82810bd0",
  2042 => x"0c81ff0b",
  2043 => x"d40c7752",
  2044 => x"87fc80d1",
  2045 => x"51bb832d",
  2046 => x"80dbc6df",
  2047 => x"5480e1b8",
  2048 => x"08802e8c",
  2049 => x"3880dbc8",
  2050 => x"5186a02d",
  2051 => x"80c0e504",
  2052 => x"81ff0bd4",
  2053 => x"0cd40870",
  2054 => x"81ff0651",
  2055 => x"537281fe",
  2056 => x"2e098106",
  2057 => x"9f3880ff",
  2058 => x"53bab42d",
  2059 => x"80e1b808",
  2060 => x"75708405",
  2061 => x"570cff13",
  2062 => x"53728025",
  2063 => x"ec388156",
  2064 => x"80c0ca04",
  2065 => x"ff145473",
  2066 => x"c73881ff",
  2067 => x"0bd40c81",
  2068 => x"ff0bd40c",
  2069 => x"d008708f",
  2070 => x"2a708106",
  2071 => x"51515372",
  2072 => x"f33872d0",
  2073 => x"0c7580e1",
  2074 => x"b80c0298",
  2075 => x"050d0402",
  2076 => x"e8050d77",
  2077 => x"797b5855",
  2078 => x"55805372",
  2079 => x"7625a538",
  2080 => x"74708105",
  2081 => x"5680f52d",
  2082 => x"74708105",
  2083 => x"5680f52d",
  2084 => x"52527171",
  2085 => x"2e873881",
  2086 => x"5180c1a6",
  2087 => x"04811353",
  2088 => x"80c0fb04",
  2089 => x"80517080",
  2090 => x"e1b80c02",
  2091 => x"98050d04",
  2092 => x"02ec050d",
  2093 => x"7680e8e4",
  2094 => x"55559f53",
  2095 => x"80747084",
  2096 => x"05560cff",
  2097 => x"13537280",
  2098 => x"25f23874",
  2099 => x"802e80c4",
  2100 => x"389a1580",
  2101 => x"e02d5180",
  2102 => x"d1c22d80",
  2103 => x"e1b80880",
  2104 => x"e1b80880",
  2105 => x"e8d80c80",
  2106 => x"e1b80854",
  2107 => x"5480e8b4",
  2108 => x"08802e9b",
  2109 => x"38941580",
  2110 => x"e02d5180",
  2111 => x"d1c22d80",
  2112 => x"e1b80890",
  2113 => x"2b83fff0",
  2114 => x"0a067075",
  2115 => x"07515372",
  2116 => x"80e8d80c",
  2117 => x"80e8d808",
  2118 => x"5372802e",
  2119 => x"9e3880e8",
  2120 => x"ac08fe14",
  2121 => x"712980e8",
  2122 => x"c0080580",
  2123 => x"e8dc0c70",
  2124 => x"842b80e8",
  2125 => x"b80c5480",
  2126 => x"c2ea0480",
  2127 => x"e8c40880",
  2128 => x"e8d80c80",
  2129 => x"e8c80880",
  2130 => x"e8dc0c80",
  2131 => x"e8b40880",
  2132 => x"2e8c3880",
  2133 => x"e8ac0884",
  2134 => x"2b5380c2",
  2135 => x"e50480e8",
  2136 => x"cc08842b",
  2137 => x"537280e8",
  2138 => x"b80c0294",
  2139 => x"050d0402",
  2140 => x"d8050d80",
  2141 => x"0b80e8b4",
  2142 => x"0c8454bc",
  2143 => x"c72d80e1",
  2144 => x"b808802e",
  2145 => x"983880e2",
  2146 => x"a8528051",
  2147 => x"bfc92d80",
  2148 => x"e1b80880",
  2149 => x"2e8738fe",
  2150 => x"5480c3a5",
  2151 => x"04ff1454",
  2152 => x"738024d7",
  2153 => x"38738e38",
  2154 => x"80dbd851",
  2155 => x"86a02d73",
  2156 => x"5580c988",
  2157 => x"04805681",
  2158 => x"0b80e8e0",
  2159 => x"0c885380",
  2160 => x"dbec5280",
  2161 => x"e2de5180",
  2162 => x"c0ef2d80",
  2163 => x"e1b80876",
  2164 => x"2e098106",
  2165 => x"893880e1",
  2166 => x"b80880e8",
  2167 => x"e00c8853",
  2168 => x"80dbf852",
  2169 => x"80e2fa51",
  2170 => x"80c0ef2d",
  2171 => x"80e1b808",
  2172 => x"893880e1",
  2173 => x"b80880e8",
  2174 => x"e00c80e8",
  2175 => x"e008802e",
  2176 => x"81843880",
  2177 => x"e5ee0b80",
  2178 => x"f52d80e5",
  2179 => x"ef0b80f5",
  2180 => x"2d71982b",
  2181 => x"71902b07",
  2182 => x"80e5f00b",
  2183 => x"80f52d70",
  2184 => x"882b7207",
  2185 => x"80e5f10b",
  2186 => x"80f52d71",
  2187 => x"0780e6a6",
  2188 => x"0b80f52d",
  2189 => x"80e6a70b",
  2190 => x"80f52d71",
  2191 => x"882b0753",
  2192 => x"5f54525a",
  2193 => x"56575573",
  2194 => x"81abaa2e",
  2195 => x"09810690",
  2196 => x"38755180",
  2197 => x"d1912d80",
  2198 => x"e1b80856",
  2199 => x"80c4ef04",
  2200 => x"7382d4d5",
  2201 => x"2e893880",
  2202 => x"dc845180",
  2203 => x"c5be0480",
  2204 => x"e2a85275",
  2205 => x"51bfc92d",
  2206 => x"80e1b808",
  2207 => x"5580e1b8",
  2208 => x"08802e84",
  2209 => x"83388853",
  2210 => x"80dbf852",
  2211 => x"80e2fa51",
  2212 => x"80c0ef2d",
  2213 => x"80e1b808",
  2214 => x"8b38810b",
  2215 => x"80e8b40c",
  2216 => x"80c5c504",
  2217 => x"885380db",
  2218 => x"ec5280e2",
  2219 => x"de5180c0",
  2220 => x"ef2d80e1",
  2221 => x"b808802e",
  2222 => x"8c3880dc",
  2223 => x"985186a0",
  2224 => x"2d80c6a4",
  2225 => x"0480e6a6",
  2226 => x"0b80f52d",
  2227 => x"547380d5",
  2228 => x"2e098106",
  2229 => x"80ce3880",
  2230 => x"e6a70b80",
  2231 => x"f52d5473",
  2232 => x"81aa2e09",
  2233 => x"8106bd38",
  2234 => x"800b80e2",
  2235 => x"a80b80f5",
  2236 => x"2d565474",
  2237 => x"81e92e83",
  2238 => x"38815474",
  2239 => x"81eb2e8c",
  2240 => x"38805573",
  2241 => x"752e0981",
  2242 => x"0682fd38",
  2243 => x"80e2b30b",
  2244 => x"80f52d55",
  2245 => x"748e3880",
  2246 => x"e2b40b80",
  2247 => x"f52d5473",
  2248 => x"822e8738",
  2249 => x"805580c9",
  2250 => x"880480e2",
  2251 => x"b50b80f5",
  2252 => x"2d7080e8",
  2253 => x"ac0cff05",
  2254 => x"80e8b00c",
  2255 => x"80e2b60b",
  2256 => x"80f52d80",
  2257 => x"e2b70b80",
  2258 => x"f52d5876",
  2259 => x"05778280",
  2260 => x"29057080",
  2261 => x"e8bc0c80",
  2262 => x"e2b80b80",
  2263 => x"f52d7080",
  2264 => x"e8d00c80",
  2265 => x"e8b40859",
  2266 => x"57587680",
  2267 => x"2e81b938",
  2268 => x"885380db",
  2269 => x"f85280e2",
  2270 => x"fa5180c0",
  2271 => x"ef2d80e1",
  2272 => x"b8088284",
  2273 => x"3880e8ac",
  2274 => x"0870842b",
  2275 => x"80e8b80c",
  2276 => x"7080e8cc",
  2277 => x"0c80e2cd",
  2278 => x"0b80f52d",
  2279 => x"80e2cc0b",
  2280 => x"80f52d71",
  2281 => x"82802905",
  2282 => x"80e2ce0b",
  2283 => x"80f52d70",
  2284 => x"84808029",
  2285 => x"1280e2cf",
  2286 => x"0b80f52d",
  2287 => x"7081800a",
  2288 => x"29127080",
  2289 => x"e8d40c80",
  2290 => x"e8d00871",
  2291 => x"2980e8bc",
  2292 => x"08057080",
  2293 => x"e8c00c80",
  2294 => x"e2d50b80",
  2295 => x"f52d80e2",
  2296 => x"d40b80f5",
  2297 => x"2d718280",
  2298 => x"290580e2",
  2299 => x"d60b80f5",
  2300 => x"2d708480",
  2301 => x"80291280",
  2302 => x"e2d70b80",
  2303 => x"f52d7098",
  2304 => x"2b81f00a",
  2305 => x"06720570",
  2306 => x"80e8c40c",
  2307 => x"fe117e29",
  2308 => x"770580e8",
  2309 => x"c80c5259",
  2310 => x"5243545e",
  2311 => x"51525952",
  2312 => x"5d575957",
  2313 => x"80c98004",
  2314 => x"80e2ba0b",
  2315 => x"80f52d80",
  2316 => x"e2b90b80",
  2317 => x"f52d7182",
  2318 => x"80290570",
  2319 => x"80e8b80c",
  2320 => x"70a02983",
  2321 => x"ff057089",
  2322 => x"2a7080e8",
  2323 => x"cc0c80e2",
  2324 => x"bf0b80f5",
  2325 => x"2d80e2be",
  2326 => x"0b80f52d",
  2327 => x"71828029",
  2328 => x"057080e8",
  2329 => x"d40c7b71",
  2330 => x"291e7080",
  2331 => x"e8c80c7d",
  2332 => x"80e8c40c",
  2333 => x"730580e8",
  2334 => x"c00c555e",
  2335 => x"51515555",
  2336 => x"805180c1",
  2337 => x"b02d8155",
  2338 => x"7480e1b8",
  2339 => x"0c02a805",
  2340 => x"0d0402ec",
  2341 => x"050d7670",
  2342 => x"872c7180",
  2343 => x"ff065556",
  2344 => x"5480e8b4",
  2345 => x"088a3873",
  2346 => x"882c7481",
  2347 => x"ff065455",
  2348 => x"80e2a852",
  2349 => x"80e8bc08",
  2350 => x"1551bfc9",
  2351 => x"2d80e1b8",
  2352 => x"085480e1",
  2353 => x"b808802e",
  2354 => x"bb3880e8",
  2355 => x"b408802e",
  2356 => x"9c387284",
  2357 => x"2980e2a8",
  2358 => x"05700852",
  2359 => x"5380d191",
  2360 => x"2d80e1b8",
  2361 => x"08f00a06",
  2362 => x"5380ca82",
  2363 => x"04721080",
  2364 => x"e2a80570",
  2365 => x"80e02d52",
  2366 => x"5380d1c2",
  2367 => x"2d80e1b8",
  2368 => x"08537254",
  2369 => x"7380e1b8",
  2370 => x"0c029405",
  2371 => x"0d0402dc",
  2372 => x"050d7a7c",
  2373 => x"59558054",
  2374 => x"77742e84",
  2375 => x"3873780c",
  2376 => x"74842c80",
  2377 => x"e8dc0805",
  2378 => x"758f0654",
  2379 => x"5972819f",
  2380 => x"3880e8b4",
  2381 => x"08802e81",
  2382 => x"8d3880e8",
  2383 => x"d8085680",
  2384 => x"e8b80875",
  2385 => x"2680f738",
  2386 => x"80e8e457",
  2387 => x"739f268f",
  2388 => x"38760853",
  2389 => x"72802e87",
  2390 => x"38725680",
  2391 => x"cb8a0475",
  2392 => x"5180c992",
  2393 => x"2d80e1b8",
  2394 => x"0880e1b8",
  2395 => x"0880ffff",
  2396 => x"fff80654",
  2397 => x"567280ff",
  2398 => x"fffff82e",
  2399 => x"83893873",
  2400 => x"9f268738",
  2401 => x"80e1b808",
  2402 => x"770c80e8",
  2403 => x"b8087571",
  2404 => x"31811684",
  2405 => x"1a5a5656",
  2406 => x"53747327",
  2407 => x"ffae3873",
  2408 => x"802e9b38",
  2409 => x"fe1680e8",
  2410 => x"ac082980",
  2411 => x"e8c00805",
  2412 => x"75842c05",
  2413 => x"7680dfd0",
  2414 => x"0c5980cb",
  2415 => x"c60480e8",
  2416 => x"d80880df",
  2417 => x"d00c80e2",
  2418 => x"a8527851",
  2419 => x"bfc92d74",
  2420 => x"852b83e0",
  2421 => x"0680e2a8",
  2422 => x"05548074",
  2423 => x"80f52d54",
  2424 => x"5672762e",
  2425 => x"09810683",
  2426 => x"38815677",
  2427 => x"802e8f38",
  2428 => x"81707706",
  2429 => x"54557280",
  2430 => x"2e843874",
  2431 => x"780c8074",
  2432 => x"80f52d56",
  2433 => x"5374732e",
  2434 => x"83388153",
  2435 => x"7481e52e",
  2436 => x"81f53881",
  2437 => x"70740654",
  2438 => x"5872802e",
  2439 => x"81e9388b",
  2440 => x"1480f52d",
  2441 => x"70832a79",
  2442 => x"06585676",
  2443 => x"9c3880df",
  2444 => x"d4085372",
  2445 => x"89387280",
  2446 => x"e6a80b81",
  2447 => x"b72d7680",
  2448 => x"dfd40c73",
  2449 => x"5380ce89",
  2450 => x"04758f2e",
  2451 => x"09810681",
  2452 => x"b638749f",
  2453 => x"068d2980",
  2454 => x"e69b1151",
  2455 => x"53811480",
  2456 => x"f52d7370",
  2457 => x"81055581",
  2458 => x"b72d8314",
  2459 => x"80f52d73",
  2460 => x"70810555",
  2461 => x"81b72d85",
  2462 => x"1480f52d",
  2463 => x"73708105",
  2464 => x"5581b72d",
  2465 => x"871480f5",
  2466 => x"2d737081",
  2467 => x"055581b7",
  2468 => x"2d891480",
  2469 => x"f52d7370",
  2470 => x"81055581",
  2471 => x"b72d8e14",
  2472 => x"80f52d73",
  2473 => x"70810555",
  2474 => x"81b72d90",
  2475 => x"1480f52d",
  2476 => x"73708105",
  2477 => x"5581b72d",
  2478 => x"921480f5",
  2479 => x"2d737081",
  2480 => x"055581b7",
  2481 => x"2d941480",
  2482 => x"f52d7370",
  2483 => x"81055581",
  2484 => x"b72d9614",
  2485 => x"80f52d73",
  2486 => x"70810555",
  2487 => x"81b72d98",
  2488 => x"1480f52d",
  2489 => x"73708105",
  2490 => x"5581b72d",
  2491 => x"9c1480f5",
  2492 => x"2d737081",
  2493 => x"055581b7",
  2494 => x"2d9e1480",
  2495 => x"f52d7381",
  2496 => x"b72d7780",
  2497 => x"dfd40c80",
  2498 => x"537280e1",
  2499 => x"b80c02a4",
  2500 => x"050d0402",
  2501 => x"cc050d7e",
  2502 => x"605e5a80",
  2503 => x"0b80e8d8",
  2504 => x"0880e8dc",
  2505 => x"08595c56",
  2506 => x"805880e8",
  2507 => x"b808782e",
  2508 => x"81bd3877",
  2509 => x"8f06a017",
  2510 => x"57547391",
  2511 => x"3880e2a8",
  2512 => x"52765181",
  2513 => x"1757bfc9",
  2514 => x"2d80e2a8",
  2515 => x"56807680",
  2516 => x"f52d5654",
  2517 => x"74742e83",
  2518 => x"38815474",
  2519 => x"81e52e81",
  2520 => x"82388170",
  2521 => x"7506555c",
  2522 => x"73802e80",
  2523 => x"f6388b16",
  2524 => x"80f52d98",
  2525 => x"06597880",
  2526 => x"ea388b53",
  2527 => x"7c527551",
  2528 => x"80c0ef2d",
  2529 => x"80e1b808",
  2530 => x"80d9389c",
  2531 => x"16085180",
  2532 => x"d1912d80",
  2533 => x"e1b80884",
  2534 => x"1b0c9a16",
  2535 => x"80e02d51",
  2536 => x"80d1c22d",
  2537 => x"80e1b808",
  2538 => x"80e1b808",
  2539 => x"881c0c80",
  2540 => x"e1b80855",
  2541 => x"5580e8b4",
  2542 => x"08802e9a",
  2543 => x"38941680",
  2544 => x"e02d5180",
  2545 => x"d1c22d80",
  2546 => x"e1b80890",
  2547 => x"2b83fff0",
  2548 => x"0a067016",
  2549 => x"51547388",
  2550 => x"1b0c787a",
  2551 => x"0c7b5480",
  2552 => x"d0ad0481",
  2553 => x"185880e8",
  2554 => x"b8087826",
  2555 => x"fec53880",
  2556 => x"e8b40880",
  2557 => x"2eb5387a",
  2558 => x"5180c992",
  2559 => x"2d80e1b8",
  2560 => x"0880e1b8",
  2561 => x"0880ffff",
  2562 => x"fff80655",
  2563 => x"5b7380ff",
  2564 => x"fffff82e",
  2565 => x"963880e1",
  2566 => x"b808fe05",
  2567 => x"80e8ac08",
  2568 => x"2980e8c0",
  2569 => x"08055780",
  2570 => x"cea80480",
  2571 => x"547380e1",
  2572 => x"b80c02b4",
  2573 => x"050d0402",
  2574 => x"f4050d74",
  2575 => x"70088105",
  2576 => x"710c7008",
  2577 => x"80e8b008",
  2578 => x"06535371",
  2579 => x"90388813",
  2580 => x"085180c9",
  2581 => x"922d80e1",
  2582 => x"b8088814",
  2583 => x"0c810b80",
  2584 => x"e1b80c02",
  2585 => x"8c050d04",
  2586 => x"02f0050d",
  2587 => x"75881108",
  2588 => x"fe0580e8",
  2589 => x"ac082980",
  2590 => x"e8c00811",
  2591 => x"720880e8",
  2592 => x"b0080605",
  2593 => x"79555354",
  2594 => x"54bfc92d",
  2595 => x"0290050d",
  2596 => x"0402f405",
  2597 => x"0d747088",
  2598 => x"2a83fe80",
  2599 => x"06707298",
  2600 => x"2a077288",
  2601 => x"2b87fc80",
  2602 => x"80067398",
  2603 => x"2b81f00a",
  2604 => x"06717307",
  2605 => x"0780e1b8",
  2606 => x"0c565153",
  2607 => x"51028c05",
  2608 => x"0d0402f8",
  2609 => x"050d028e",
  2610 => x"0580f52d",
  2611 => x"74882b07",
  2612 => x"7083ffff",
  2613 => x"0680e1b8",
  2614 => x"0c510288",
  2615 => x"050d0402",
  2616 => x"f4050d74",
  2617 => x"76785354",
  2618 => x"52807125",
  2619 => x"97387270",
  2620 => x"81055480",
  2621 => x"f52d7270",
  2622 => x"81055481",
  2623 => x"b72dff11",
  2624 => x"5170eb38",
  2625 => x"807281b7",
  2626 => x"2d028c05",
  2627 => x"0d0402e0",
  2628 => x"050d7957",
  2629 => x"80705970",
  2630 => x"575580d2",
  2631 => x"c50402a0",
  2632 => x"05fc0552",
  2633 => x"755180ca",
  2634 => x"8e2d80e1",
  2635 => x"b80880e1",
  2636 => x"b8080981",
  2637 => x"057080e1",
  2638 => x"b808079f",
  2639 => x"2a770581",
  2640 => x"19595754",
  2641 => x"54767525",
  2642 => x"53778438",
  2643 => x"72d03873",
  2644 => x"80e1b80c",
  2645 => x"02a0050d",
  2646 => x"0402f005",
  2647 => x"0d80e1b4",
  2648 => x"08165180",
  2649 => x"d28e2d80",
  2650 => x"e1b80880",
  2651 => x"2ea0388b",
  2652 => x"5380e1b8",
  2653 => x"085280e6",
  2654 => x"a85180d1",
  2655 => x"df2d80e9",
  2656 => x"e4085473",
  2657 => x"802e8738",
  2658 => x"80e6a851",
  2659 => x"732d0290",
  2660 => x"050d0402",
  2661 => x"f4050d74",
  2662 => x"76708c2c",
  2663 => x"708f0680",
  2664 => x"dcc80805",
  2665 => x"51535353",
  2666 => x"7080f52d",
  2667 => x"7381b72d",
  2668 => x"71882c70",
  2669 => x"8f0680dc",
  2670 => x"c8080551",
  2671 => x"517080f5",
  2672 => x"2d811481",
  2673 => x"b72d7184",
  2674 => x"2c708f06",
  2675 => x"80dcc808",
  2676 => x"05515170",
  2677 => x"80f52d82",
  2678 => x"1481b72d",
  2679 => x"718f0680",
  2680 => x"dcc80805",
  2681 => x"527180f5",
  2682 => x"2d831481",
  2683 => x"b72d028c",
  2684 => x"050d0402",
  2685 => x"d8050d80",
  2686 => x"5a807056",
  2687 => x"5980d4a3",
  2688 => x"0402a805",
  2689 => x"fc055278",
  2690 => x"5180ca8e",
  2691 => x"2d80e1b8",
  2692 => x"08098105",
  2693 => x"7080e1b8",
  2694 => x"08079f2a",
  2695 => x"7605811b",
  2696 => x"5b565480",
  2697 => x"e1b40875",
  2698 => x"24547984",
  2699 => x"3873d238",
  2700 => x"80705b55",
  2701 => x"02a805fc",
  2702 => x"05527851",
  2703 => x"80ca8e2d",
  2704 => x"80e1b808",
  2705 => x"802e81b4",
  2706 => x"3880e1b8",
  2707 => x"088b0580",
  2708 => x"f52d7084",
  2709 => x"2a708106",
  2710 => x"77107884",
  2711 => x"2b80e6a8",
  2712 => x"0b80f52d",
  2713 => x"5c5c5351",
  2714 => x"55567380",
  2715 => x"2e80ce38",
  2716 => x"7416822b",
  2717 => x"80d8920b",
  2718 => x"80dfe012",
  2719 => x"0c547775",
  2720 => x"311080e9",
  2721 => x"e8115556",
  2722 => x"90747081",
  2723 => x"055681b7",
  2724 => x"2da07481",
  2725 => x"b72d7681",
  2726 => x"ff068116",
  2727 => x"58547380",
  2728 => x"2e8b389c",
  2729 => x"5380e6a8",
  2730 => x"5280d5b4",
  2731 => x"048b5380",
  2732 => x"e1b80852",
  2733 => x"80e9ea16",
  2734 => x"5180d5f2",
  2735 => x"04741682",
  2736 => x"2b80d2d9",
  2737 => x"0b80dfe0",
  2738 => x"120c5476",
  2739 => x"81ff0681",
  2740 => x"16585473",
  2741 => x"802e8b38",
  2742 => x"9c5380e6",
  2743 => x"a85280d5",
  2744 => x"e9048b53",
  2745 => x"80e1b808",
  2746 => x"52777531",
  2747 => x"1080e9e8",
  2748 => x"05517655",
  2749 => x"80d1df2d",
  2750 => x"80d69104",
  2751 => x"74902975",
  2752 => x"31701080",
  2753 => x"e9e80551",
  2754 => x"5480e1b8",
  2755 => x"087481b7",
  2756 => x"2d811959",
  2757 => x"748b24a6",
  2758 => x"3879802e",
  2759 => x"fe963874",
  2760 => x"90297531",
  2761 => x"701080e9",
  2762 => x"e8058c77",
  2763 => x"31575154",
  2764 => x"807481b7",
  2765 => x"2d9e14ff",
  2766 => x"16565474",
  2767 => x"f33880dc",
  2768 => x"a45280e1",
  2769 => x"8c51a290",
  2770 => x"2d80e1b4",
  2771 => x"085280e1",
  2772 => x"915180d3",
  2773 => x"932d80e8",
  2774 => x"b8085280",
  2775 => x"e1965180",
  2776 => x"d3932d78",
  2777 => x"5280e19b",
  2778 => x"5180d393",
  2779 => x"2d80dfd0",
  2780 => x"0b80e02d",
  2781 => x"5280e1a0",
  2782 => x"5180d393",
  2783 => x"2d80dfd2",
  2784 => x"0b80e02d",
  2785 => x"5280e1a4",
  2786 => x"5180d393",
  2787 => x"2d7880e1",
  2788 => x"b80c02a8",
  2789 => x"050d0402",
  2790 => x"fc050d72",
  2791 => x"5170fd2e",
  2792 => x"b23870fd",
  2793 => x"248b3870",
  2794 => x"fc2e80d0",
  2795 => x"3880d886",
  2796 => x"0470fe2e",
  2797 => x"b93870ff",
  2798 => x"2e098106",
  2799 => x"80c83880",
  2800 => x"e1b40851",
  2801 => x"70802ebe",
  2802 => x"38ff1180",
  2803 => x"e1b40c80",
  2804 => x"d8860480",
  2805 => x"e1b408f4",
  2806 => x"057080e1",
  2807 => x"b40c5170",
  2808 => x"8025a338",
  2809 => x"800b80e1",
  2810 => x"b40c80d8",
  2811 => x"860480e1",
  2812 => x"b4088105",
  2813 => x"80e1b40c",
  2814 => x"80d88604",
  2815 => x"80e1b408",
  2816 => x"8c0580e1",
  2817 => x"b40c80d3",
  2818 => x"f32dafb6",
  2819 => x"2d028405",
  2820 => x"0d0402fc",
  2821 => x"050d80e1",
  2822 => x"b4081351",
  2823 => x"80d28e2d",
  2824 => x"80e1b808",
  2825 => x"802e8a38",
  2826 => x"80e1b808",
  2827 => x"5180c1b0",
  2828 => x"2d800b80",
  2829 => x"e1b40c80",
  2830 => x"d3f32daf",
  2831 => x"b62d0284",
  2832 => x"050d0402",
  2833 => x"fc050d80",
  2834 => x"0b80e1b4",
  2835 => x"0c80d3f3",
  2836 => x"2daeb22d",
  2837 => x"80e1b808",
  2838 => x"80e0fc0c",
  2839 => x"80dfd851",
  2840 => x"b0dc2d02",
  2841 => x"84050d04",
  2842 => x"7180e9e4",
  2843 => x"0c040000",
  2844 => x"00ffffff",
  2845 => x"ff00ffff",
  2846 => x"ffff00ff",
  2847 => x"ffffff00",
  2848 => x"30313233",
  2849 => x"34353637",
  2850 => x"38394142",
  2851 => x"43444546",
  2852 => x"00000000",
  2853 => x"52657365",
  2854 => x"74000000",
  2855 => x"5363616e",
  2856 => x"6c696e65",
  2857 => x"73000000",
  2858 => x"50414c20",
  2859 => x"2f204e54",
  2860 => x"53430000",
  2861 => x"436f6c6f",
  2862 => x"72000000",
  2863 => x"44696666",
  2864 => x"6963756c",
  2865 => x"74792041",
  2866 => x"00000000",
  2867 => x"44696666",
  2868 => x"6963756c",
  2869 => x"74792042",
  2870 => x"00000000",
  2871 => x"2a537570",
  2872 => x"65726368",
  2873 => x"69702069",
  2874 => x"6e206361",
  2875 => x"72747269",
  2876 => x"64676500",
  2877 => x"2a42616e",
  2878 => x"6b204530",
  2879 => x"00000000",
  2880 => x"2a42616e",
  2881 => x"6b204537",
  2882 => x"00000000",
  2883 => x"53656c65",
  2884 => x"63740000",
  2885 => x"53746172",
  2886 => x"74000000",
  2887 => x"4c6f6164",
  2888 => x"20524f4d",
  2889 => x"20100000",
  2890 => x"45786974",
  2891 => x"00000000",
  2892 => x"524f4d20",
  2893 => x"6c6f6164",
  2894 => x"696e6720",
  2895 => x"6661696c",
  2896 => x"65640000",
  2897 => x"4f4b0000",
  2898 => x"496e6974",
  2899 => x"69616c69",
  2900 => x"7a696e67",
  2901 => x"20534420",
  2902 => x"63617264",
  2903 => x"0a000000",
  2904 => x"446f6e65",
  2905 => x"20696e69",
  2906 => x"7469616c",
  2907 => x"697a6174",
  2908 => x"696f6e0a",
  2909 => x"00000000",
  2910 => x"16200000",
  2911 => x"14200000",
  2912 => x"15200000",
  2913 => x"53442069",
  2914 => x"6e69742e",
  2915 => x"2e2e0a00",
  2916 => x"53442063",
  2917 => x"61726420",
  2918 => x"72657365",
  2919 => x"74206661",
  2920 => x"696c6564",
  2921 => x"210a0000",
  2922 => x"53444843",
  2923 => x"20657272",
  2924 => x"6f72210a",
  2925 => x"00000000",
  2926 => x"57726974",
  2927 => x"65206661",
  2928 => x"696c6564",
  2929 => x"0a000000",
  2930 => x"52656164",
  2931 => x"20666169",
  2932 => x"6c65640a",
  2933 => x"00000000",
  2934 => x"43617264",
  2935 => x"20696e69",
  2936 => x"74206661",
  2937 => x"696c6564",
  2938 => x"0a000000",
  2939 => x"46415431",
  2940 => x"36202020",
  2941 => x"00000000",
  2942 => x"46415433",
  2943 => x"32202020",
  2944 => x"00000000",
  2945 => x"4e6f2070",
  2946 => x"61727469",
  2947 => x"74696f6e",
  2948 => x"20736967",
  2949 => x"0a000000",
  2950 => x"42616420",
  2951 => x"70617274",
  2952 => x"0a000000",
  2953 => x"4261636b",
  2954 => x"20787878",
  2955 => x"78207979",
  2956 => x"7979207a",
  2957 => x"7a7a7a20",
  2958 => x"6b6b6b6b",
  2959 => x"6b6b6b6b",
  2960 => x"00000000",
  2961 => x"00000002",
  2962 => x"00002c80",
  2963 => x"00000002",
  2964 => x"00002c94",
  2965 => x"0000035a",
  2966 => x"00000001",
  2967 => x"00002c9c",
  2968 => x"00000000",
  2969 => x"00000001",
  2970 => x"00002ca8",
  2971 => x"00000001",
  2972 => x"00000001",
  2973 => x"00002cb4",
  2974 => x"00000002",
  2975 => x"00000001",
  2976 => x"00002cbc",
  2977 => x"00000003",
  2978 => x"00000001",
  2979 => x"00002ccc",
  2980 => x"00000004",
  2981 => x"00000001",
  2982 => x"00002cdc",
  2983 => x"00000005",
  2984 => x"00000001",
  2985 => x"00002cf4",
  2986 => x"00000008",
  2987 => x"00000001",
  2988 => x"00002d00",
  2989 => x"00000009",
  2990 => x"00000002",
  2991 => x"00002d0c",
  2992 => x"0000036e",
  2993 => x"00000002",
  2994 => x"00002d14",
  2995 => x"00000a3f",
  2996 => x"00000002",
  2997 => x"00002d1c",
  2998 => x"00002c43",
  2999 => x"00000002",
  3000 => x"00002d28",
  3001 => x"0000174f",
  3002 => x"00000000",
  3003 => x"00000000",
  3004 => x"00000000",
  3005 => x"00000004",
  3006 => x"00002d30",
  3007 => x"00002ef4",
  3008 => x"00000004",
  3009 => x"00002d44",
  3010 => x"00002e4c",
  3011 => x"00000000",
  3012 => x"00000000",
  3013 => x"00000000",
  3014 => x"00000000",
  3015 => x"00000000",
  3016 => x"00000000",
  3017 => x"00000000",
  3018 => x"00000000",
  3019 => x"00000000",
  3020 => x"00000000",
  3021 => x"00000000",
  3022 => x"00000000",
  3023 => x"00000000",
  3024 => x"00000000",
  3025 => x"00000000",
  3026 => x"00000000",
  3027 => x"00000000",
  3028 => x"00000000",
  3029 => x"00000000",
  3030 => x"761c1c1c",
  3031 => x"1c1c051c",
  3032 => x"1c1c1c1c",
  3033 => x"f2f5fafd",
  3034 => x"5a000000",
  3035 => x"00000000",
  3036 => x"00000000",
  3037 => x"00000000",
  3038 => x"00000000",
  3039 => x"00000000",
  3040 => x"00000000",
  3041 => x"00000000",
  3042 => x"00000000",
  3043 => x"00000000",
  3044 => x"00000000",
  3045 => x"00000000",
  3046 => x"00000000",
  3047 => x"00000000",
  3048 => x"00000000",
  3049 => x"00000000",
  3050 => x"00000000",
  3051 => x"00000000",
  3052 => x"00000000",
  3053 => x"0001ffff",
  3054 => x"0001ffff",
  3055 => x"0001ffff",
  3056 => x"00000000",
  3057 => x"00000000",
  3058 => x"00000004",
  3059 => x"00000000",
  3060 => x"00000000",
  3061 => x"00000000",
  3062 => x"00000002",
  3063 => x"000034e8",
  3064 => x"00002959",
  3065 => x"00000002",
  3066 => x"00003506",
  3067 => x"00002959",
  3068 => x"00000002",
  3069 => x"00003524",
  3070 => x"00002959",
  3071 => x"00000002",
  3072 => x"00003542",
  3073 => x"00002959",
  3074 => x"00000002",
  3075 => x"00003560",
  3076 => x"00002959",
  3077 => x"00000002",
  3078 => x"0000357e",
  3079 => x"00002959",
  3080 => x"00000002",
  3081 => x"0000359c",
  3082 => x"00002959",
  3083 => x"00000002",
  3084 => x"000035ba",
  3085 => x"00002959",
  3086 => x"00000002",
  3087 => x"000035d8",
  3088 => x"00002959",
  3089 => x"00000002",
  3090 => x"000035f6",
  3091 => x"00002959",
  3092 => x"00000002",
  3093 => x"00003614",
  3094 => x"00002959",
  3095 => x"00000002",
  3096 => x"00003632",
  3097 => x"00002959",
  3098 => x"00000002",
  3099 => x"00003650",
  3100 => x"00002959",
  3101 => x"00000004",
  3102 => x"0000308c",
  3103 => x"00000000",
  3104 => x"00000000",
  3105 => x"00000000",
  3106 => x"00002b97",
  3107 => x"4261636b",
  3108 => x"00000000",
  3109 => x"00000000",
  3110 => x"00000000",
  3111 => x"00000000",
  3112 => x"00000000",
  3113 => x"00000000",
  3114 => x"00000000",
  3115 => x"00000000",
  3116 => x"00000000",
  3117 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

