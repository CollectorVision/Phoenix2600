-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80e1",
     9 => x"84080b0b",
    10 => x"80e18808",
    11 => x"0b0b80e1",
    12 => x"8c080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"e18c0c0b",
    16 => x"0b80e188",
    17 => x"0c0b0b80",
    18 => x"e1840c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d8bc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80e18470",
    57 => x"80ebbc27",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a6d9",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80e1",
    65 => x"940c9f0b",
    66 => x"80e1980c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"e19808ff",
    70 => x"0580e198",
    71 => x"0c80e198",
    72 => x"088025e8",
    73 => x"3880e194",
    74 => x"08ff0580",
    75 => x"e1940c80",
    76 => x"e1940880",
    77 => x"25d03880",
    78 => x"0b80e198",
    79 => x"0c800b80",
    80 => x"e1940c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80e19408",
   100 => x"25913882",
   101 => x"c82d80e1",
   102 => x"9408ff05",
   103 => x"80e1940c",
   104 => x"838a0480",
   105 => x"e1940880",
   106 => x"e1980853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80e19408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"e1980881",
   116 => x"0580e198",
   117 => x"0c80e198",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80e198",
   121 => x"0c80e194",
   122 => x"08810580",
   123 => x"e1940c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480e1",
   128 => x"98088105",
   129 => x"80e1980c",
   130 => x"80e19808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80e198",
   134 => x"0c80e194",
   135 => x"08810580",
   136 => x"e1940c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"e19c0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"e19c0c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280e1",
   177 => x"9c088407",
   178 => x"80e19c0c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80dc",
   183 => x"900c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80e19c",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80e1",
   208 => x"840c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02f4050d",
  1093 => x"74765452",
  1094 => x"72708105",
  1095 => x"5480f52d",
  1096 => x"51707270",
  1097 => x"81055481",
  1098 => x"b72d70ec",
  1099 => x"38707281",
  1100 => x"b72d028c",
  1101 => x"050d0402",
  1102 => x"f4050d80",
  1103 => x"dcac0b80",
  1104 => x"f52d80df",
  1105 => x"94087081",
  1106 => x"06535452",
  1107 => x"70802e85",
  1108 => x"38718407",
  1109 => x"5272812a",
  1110 => x"70810651",
  1111 => x"5170802e",
  1112 => x"85387182",
  1113 => x"07527282",
  1114 => x"2a708106",
  1115 => x"51517080",
  1116 => x"2e853871",
  1117 => x"81075272",
  1118 => x"832a7081",
  1119 => x"06515170",
  1120 => x"802e8538",
  1121 => x"71880752",
  1122 => x"72842a70",
  1123 => x"81065151",
  1124 => x"70802e85",
  1125 => x"38719007",
  1126 => x"5272852a",
  1127 => x"70810651",
  1128 => x"5170802e",
  1129 => x"853871a0",
  1130 => x"07527288",
  1131 => x"2a708106",
  1132 => x"51517080",
  1133 => x"2e863871",
  1134 => x"80c00752",
  1135 => x"72892a70",
  1136 => x"81065151",
  1137 => x"70802e86",
  1138 => x"38718180",
  1139 => x"075271fc",
  1140 => x"0c7180e1",
  1141 => x"840c028c",
  1142 => x"050d0402",
  1143 => x"cc050d7e",
  1144 => x"5d800b80",
  1145 => x"df940881",
  1146 => x"8006715c",
  1147 => x"5d5b810b",
  1148 => x"ec0c840b",
  1149 => x"ec0c7c52",
  1150 => x"80e1a051",
  1151 => x"80cddf2d",
  1152 => x"80e18408",
  1153 => x"7b2e80ff",
  1154 => x"3880e1a4",
  1155 => x"087bff12",
  1156 => x"57595774",
  1157 => x"7b2e8b38",
  1158 => x"81187581",
  1159 => x"2a565874",
  1160 => x"f738f718",
  1161 => x"58815b80",
  1162 => x"772580db",
  1163 => x"38775274",
  1164 => x"5184a82d",
  1165 => x"80e1f452",
  1166 => x"80e1a051",
  1167 => x"80d0b42d",
  1168 => x"80e18408",
  1169 => x"802ea638",
  1170 => x"80e1f459",
  1171 => x"7ba73883",
  1172 => x"ff567870",
  1173 => x"81055a80",
  1174 => x"f52d7a81",
  1175 => x"1c5ce40c",
  1176 => x"e80cff16",
  1177 => x"56758025",
  1178 => x"e938a4f5",
  1179 => x"0480e184",
  1180 => x"085b8480",
  1181 => x"5780e1a0",
  1182 => x"5180d083",
  1183 => x"2dfc8017",
  1184 => x"81165657",
  1185 => x"a4a70480",
  1186 => x"e1a408f8",
  1187 => x"0c881d54",
  1188 => x"807480f5",
  1189 => x"2d7081ff",
  1190 => x"06555855",
  1191 => x"72752eb6",
  1192 => x"38811480",
  1193 => x"f52d5372",
  1194 => x"752eab38",
  1195 => x"74821580",
  1196 => x"f52d5456",
  1197 => x"7280d32e",
  1198 => x"09810683",
  1199 => x"38815672",
  1200 => x"80f33270",
  1201 => x"09810570",
  1202 => x"80257807",
  1203 => x"51515372",
  1204 => x"802e8338",
  1205 => x"a0558077",
  1206 => x"81ff0654",
  1207 => x"567280c5",
  1208 => x"2e098106",
  1209 => x"83388156",
  1210 => x"7280e532",
  1211 => x"70098105",
  1212 => x"70802578",
  1213 => x"07515153",
  1214 => x"72802ea4",
  1215 => x"38811480",
  1216 => x"f52d5372",
  1217 => x"b02e0981",
  1218 => x"06893874",
  1219 => x"82800755",
  1220 => x"a6a00472",
  1221 => x"b72e0981",
  1222 => x"06863874",
  1223 => x"84800755",
  1224 => x"80df9408",
  1225 => x"f9df0675",
  1226 => x"0780df94",
  1227 => x"0ca2b72d",
  1228 => x"800be00c",
  1229 => x"805186da",
  1230 => x"2d86c72d",
  1231 => x"7a802e88",
  1232 => x"3880dc98",
  1233 => x"51a6cc04",
  1234 => x"80ddc051",
  1235 => x"b0dc2d7a",
  1236 => x"80e1840c",
  1237 => x"02b4050d",
  1238 => x"0402f405",
  1239 => x"0d840bec",
  1240 => x"0c810be0",
  1241 => x"0cae992d",
  1242 => x"a7f32d81",
  1243 => x"f92d8352",
  1244 => x"adfc2d81",
  1245 => x"51858d2d",
  1246 => x"ff125271",
  1247 => x"8025f138",
  1248 => x"840bec0c",
  1249 => x"80da9451",
  1250 => x"86a02d80",
  1251 => x"c2da2d80",
  1252 => x"e1840880",
  1253 => x"2e80c538",
  1254 => x"80daac51",
  1255 => x"86a02da3",
  1256 => x"db5180d8",
  1257 => x"b42d80dc",
  1258 => x"9851b0dc",
  1259 => x"2daebb2d",
  1260 => x"a99e2d80",
  1261 => x"e1840881",
  1262 => x"06527180",
  1263 => x"2e863880",
  1264 => x"5194bf2d",
  1265 => x"b0ef2d80",
  1266 => x"e1840852",
  1267 => x"a2b72d86",
  1268 => x"53718338",
  1269 => x"845372ec",
  1270 => x"0ca7b004",
  1271 => x"800b80e1",
  1272 => x"840c028c",
  1273 => x"050d0471",
  1274 => x"980c04ff",
  1275 => x"b00880e1",
  1276 => x"840c0481",
  1277 => x"0bffb00c",
  1278 => x"04800bff",
  1279 => x"b00c0402",
  1280 => x"d8050dff",
  1281 => x"b40887ff",
  1282 => x"ff065a81",
  1283 => x"54807080",
  1284 => x"df800880",
  1285 => x"df840880",
  1286 => x"dedc5b59",
  1287 => x"575a5879",
  1288 => x"74067575",
  1289 => x"06525271",
  1290 => x"712e8d38",
  1291 => x"8077818a",
  1292 => x"2d730975",
  1293 => x"06720755",
  1294 => x"7680e02d",
  1295 => x"7083ffff",
  1296 => x"06535171",
  1297 => x"80e42e09",
  1298 => x"8106a238",
  1299 => x"74740670",
  1300 => x"77760632",
  1301 => x"70098105",
  1302 => x"7072079f",
  1303 => x"2a7b0577",
  1304 => x"097a0674",
  1305 => x"075a5b53",
  1306 => x"5353a8fb",
  1307 => x"047180e4",
  1308 => x"26893881",
  1309 => x"11517077",
  1310 => x"818a2d73",
  1311 => x"10811a82",
  1312 => x"19595a54",
  1313 => x"907925ff",
  1314 => x"96387580",
  1315 => x"df840c74",
  1316 => x"80df800c",
  1317 => x"7780e184",
  1318 => x"0c02a805",
  1319 => x"0d0402d0",
  1320 => x"050d805c",
  1321 => x"aaae0480",
  1322 => x"e1840881",
  1323 => x"f02e0981",
  1324 => x"068a3881",
  1325 => x"0b80df8c",
  1326 => x"0caaae04",
  1327 => x"80e18408",
  1328 => x"81e02e09",
  1329 => x"81068a38",
  1330 => x"810b80df",
  1331 => x"900caaae",
  1332 => x"0480e184",
  1333 => x"085280df",
  1334 => x"9008802e",
  1335 => x"893880e1",
  1336 => x"84088180",
  1337 => x"05527184",
  1338 => x"2c728f06",
  1339 => x"535380df",
  1340 => x"8c08802e",
  1341 => x"9a387284",
  1342 => x"2980dde4",
  1343 => x"05721381",
  1344 => x"712b7009",
  1345 => x"73080673",
  1346 => x"0c515353",
  1347 => x"aaa20472",
  1348 => x"842980dd",
  1349 => x"e4057213",
  1350 => x"83712b72",
  1351 => x"0807720c",
  1352 => x"5353800b",
  1353 => x"80df900c",
  1354 => x"800b80df",
  1355 => x"8c0c80e1",
  1356 => x"ac51acef",
  1357 => x"2d80e184",
  1358 => x"08ff24fe",
  1359 => x"ea38a7ff",
  1360 => x"2d80e184",
  1361 => x"08802e81",
  1362 => x"b0388159",
  1363 => x"800b80df",
  1364 => x"880880df",
  1365 => x"840880de",
  1366 => x"b85a5c5c",
  1367 => x"587a7906",
  1368 => x"7a7a0654",
  1369 => x"5271732e",
  1370 => x"80f83872",
  1371 => x"09810570",
  1372 => x"74078025",
  1373 => x"80dea41a",
  1374 => x"80f52d70",
  1375 => x"842c718f",
  1376 => x"06585357",
  1377 => x"57527580",
  1378 => x"2ea33871",
  1379 => x"842980dd",
  1380 => x"e4057415",
  1381 => x"83712b72",
  1382 => x"0807720c",
  1383 => x"54527680",
  1384 => x"e02d8105",
  1385 => x"52717781",
  1386 => x"8a2dabc3",
  1387 => x"04718429",
  1388 => x"80dde405",
  1389 => x"74158171",
  1390 => x"2b700973",
  1391 => x"0806730c",
  1392 => x"51535374",
  1393 => x"85327009",
  1394 => x"81057080",
  1395 => x"25515152",
  1396 => x"75802e8e",
  1397 => x"38817073",
  1398 => x"06535371",
  1399 => x"802e8338",
  1400 => x"725c7810",
  1401 => x"81198219",
  1402 => x"59595990",
  1403 => x"7825feed",
  1404 => x"3880df84",
  1405 => x"0880df88",
  1406 => x"0c7b80e1",
  1407 => x"840c02b0",
  1408 => x"050d0402",
  1409 => x"f8050d80",
  1410 => x"dde4528f",
  1411 => x"51807270",
  1412 => x"8405540c",
  1413 => x"ff115170",
  1414 => x"8025f238",
  1415 => x"0288050d",
  1416 => x"0402f005",
  1417 => x"0d7551a7",
  1418 => x"f92d7082",
  1419 => x"2cfc0680",
  1420 => x"dde41172",
  1421 => x"109e0671",
  1422 => x"0870722a",
  1423 => x"70830682",
  1424 => x"742b7009",
  1425 => x"7406760c",
  1426 => x"54515657",
  1427 => x"535153a7",
  1428 => x"f32d7180",
  1429 => x"e1840c02",
  1430 => x"90050d04",
  1431 => x"02fc050d",
  1432 => x"72518071",
  1433 => x"0c800b84",
  1434 => x"120c0284",
  1435 => x"050d0402",
  1436 => x"f0050d75",
  1437 => x"70088412",
  1438 => x"08535353",
  1439 => x"ff547171",
  1440 => x"2ea838a7",
  1441 => x"f92d8413",
  1442 => x"08708429",
  1443 => x"14881170",
  1444 => x"087081ff",
  1445 => x"06841808",
  1446 => x"81118706",
  1447 => x"841a0c53",
  1448 => x"51555151",
  1449 => x"51a7f32d",
  1450 => x"71547380",
  1451 => x"e1840c02",
  1452 => x"90050d04",
  1453 => x"02f8050d",
  1454 => x"a7f92de0",
  1455 => x"08708b2a",
  1456 => x"70810651",
  1457 => x"52527080",
  1458 => x"2ea13880",
  1459 => x"e1ac0870",
  1460 => x"842980e1",
  1461 => x"b4057381",
  1462 => x"ff06710c",
  1463 => x"515180e1",
  1464 => x"ac088111",
  1465 => x"870680e1",
  1466 => x"ac0c5180",
  1467 => x"0b80e1d4",
  1468 => x"0ca7eb2d",
  1469 => x"a7f32d02",
  1470 => x"88050d04",
  1471 => x"02fc050d",
  1472 => x"a7f92d81",
  1473 => x"0b80e1d4",
  1474 => x"0ca7f32d",
  1475 => x"80e1d408",
  1476 => x"5170f938",
  1477 => x"0284050d",
  1478 => x"0402fc05",
  1479 => x"0d80e1ac",
  1480 => x"51acdc2d",
  1481 => x"ac832dad",
  1482 => x"b451a7e7",
  1483 => x"2d028405",
  1484 => x"0d0480e1",
  1485 => x"e00880e1",
  1486 => x"840c0402",
  1487 => x"fc050d81",
  1488 => x"0b80df98",
  1489 => x"0c815185",
  1490 => x"8d2d0284",
  1491 => x"050d0402",
  1492 => x"fc050dae",
  1493 => x"d904a99e",
  1494 => x"2d80f651",
  1495 => x"aca12d80",
  1496 => x"e18408f2",
  1497 => x"3880da51",
  1498 => x"aca12d80",
  1499 => x"e18408e6",
  1500 => x"3880e184",
  1501 => x"0880df98",
  1502 => x"0c80e184",
  1503 => x"0851858d",
  1504 => x"2d028405",
  1505 => x"0d0402ec",
  1506 => x"050d7654",
  1507 => x"8052870b",
  1508 => x"881580f5",
  1509 => x"2d565374",
  1510 => x"72248338",
  1511 => x"a0537251",
  1512 => x"83842d81",
  1513 => x"128b1580",
  1514 => x"f52d5452",
  1515 => x"727225de",
  1516 => x"38029405",
  1517 => x"0d0402f0",
  1518 => x"050d80e1",
  1519 => x"e0085481",
  1520 => x"f92d800b",
  1521 => x"80e1e40c",
  1522 => x"7308802e",
  1523 => x"81893882",
  1524 => x"0b80e198",
  1525 => x"0c80e1e4",
  1526 => x"088f0680",
  1527 => x"e1940c73",
  1528 => x"08527183",
  1529 => x"2e963871",
  1530 => x"83268938",
  1531 => x"71812eb0",
  1532 => x"38b0c004",
  1533 => x"71852ea0",
  1534 => x"38b0c004",
  1535 => x"881480f5",
  1536 => x"2d841508",
  1537 => x"80dac453",
  1538 => x"545286a0",
  1539 => x"2d718429",
  1540 => x"13700852",
  1541 => x"52b0c404",
  1542 => x"7351af86",
  1543 => x"2db0c004",
  1544 => x"80df9408",
  1545 => x"8815082c",
  1546 => x"70810651",
  1547 => x"5271802e",
  1548 => x"883880da",
  1549 => x"c851b0bd",
  1550 => x"0480dacc",
  1551 => x"5186a02d",
  1552 => x"84140851",
  1553 => x"86a02d80",
  1554 => x"e1e40881",
  1555 => x"0580e1e4",
  1556 => x"0c8c1454",
  1557 => x"afc80402",
  1558 => x"90050d04",
  1559 => x"7180e1e0",
  1560 => x"0cafb62d",
  1561 => x"80e1e408",
  1562 => x"ff0580e1",
  1563 => x"e80c0402",
  1564 => x"e8050d80",
  1565 => x"e1e00880",
  1566 => x"e1ec0857",
  1567 => x"5580f651",
  1568 => x"aca12d80",
  1569 => x"e1840881",
  1570 => x"2a708106",
  1571 => x"51527180",
  1572 => x"2ea438b1",
  1573 => x"9904a99e",
  1574 => x"2d80f651",
  1575 => x"aca12d80",
  1576 => x"e18408f2",
  1577 => x"3880df98",
  1578 => x"08813270",
  1579 => x"80df980c",
  1580 => x"70525285",
  1581 => x"8d2d800b",
  1582 => x"80e1d80c",
  1583 => x"800b80e1",
  1584 => x"dc0c80df",
  1585 => x"9808838d",
  1586 => x"3880da51",
  1587 => x"aca12d80",
  1588 => x"e1840880",
  1589 => x"2e8c3880",
  1590 => x"e1d80881",
  1591 => x"800780e1",
  1592 => x"d80c80d9",
  1593 => x"51aca12d",
  1594 => x"80e18408",
  1595 => x"802e8c38",
  1596 => x"80e1d808",
  1597 => x"80c00780",
  1598 => x"e1d80c81",
  1599 => x"9451aca1",
  1600 => x"2d80e184",
  1601 => x"08802e8b",
  1602 => x"3880e1d8",
  1603 => x"08900780",
  1604 => x"e1d80c81",
  1605 => x"9151aca1",
  1606 => x"2d80e184",
  1607 => x"08802e8b",
  1608 => x"3880e1d8",
  1609 => x"08a00780",
  1610 => x"e1d80c81",
  1611 => x"f551aca1",
  1612 => x"2d80e184",
  1613 => x"08802e8b",
  1614 => x"3880e1d8",
  1615 => x"08810780",
  1616 => x"e1d80c81",
  1617 => x"f251aca1",
  1618 => x"2d80e184",
  1619 => x"08802e8b",
  1620 => x"3880e1d8",
  1621 => x"08820780",
  1622 => x"e1d80c81",
  1623 => x"eb51aca1",
  1624 => x"2d80e184",
  1625 => x"08802e8b",
  1626 => x"3880e1d8",
  1627 => x"08840780",
  1628 => x"e1d80c81",
  1629 => x"f451aca1",
  1630 => x"2d80e184",
  1631 => x"08802e8b",
  1632 => x"3880e1d8",
  1633 => x"08880780",
  1634 => x"e1d80c80",
  1635 => x"d851aca1",
  1636 => x"2d80e184",
  1637 => x"08802e8c",
  1638 => x"3880e1dc",
  1639 => x"08818007",
  1640 => x"80e1dc0c",
  1641 => x"9251aca1",
  1642 => x"2d80e184",
  1643 => x"08802e8c",
  1644 => x"3880e1dc",
  1645 => x"0880c007",
  1646 => x"80e1dc0c",
  1647 => x"9451aca1",
  1648 => x"2d80e184",
  1649 => x"08802e8b",
  1650 => x"3880e1dc",
  1651 => x"08900780",
  1652 => x"e1dc0c91",
  1653 => x"51aca12d",
  1654 => x"80e18408",
  1655 => x"802e8b38",
  1656 => x"80e1dc08",
  1657 => x"a00780e1",
  1658 => x"dc0c9d51",
  1659 => x"aca12d80",
  1660 => x"e1840880",
  1661 => x"2e8b3880",
  1662 => x"e1dc0881",
  1663 => x"0780e1dc",
  1664 => x"0c9b51ac",
  1665 => x"a12d80e1",
  1666 => x"8408802e",
  1667 => x"8b3880e1",
  1668 => x"dc088207",
  1669 => x"80e1dc0c",
  1670 => x"9c51aca1",
  1671 => x"2d80e184",
  1672 => x"08802e8b",
  1673 => x"3880e1dc",
  1674 => x"08840780",
  1675 => x"e1dc0ca3",
  1676 => x"51aca12d",
  1677 => x"80e18408",
  1678 => x"802e8b38",
  1679 => x"80e1dc08",
  1680 => x"880780e1",
  1681 => x"dc0c81fd",
  1682 => x"51aca12d",
  1683 => x"81fa51ac",
  1684 => x"a12dbaaa",
  1685 => x"0481f551",
  1686 => x"aca12d80",
  1687 => x"e1840881",
  1688 => x"2a708106",
  1689 => x"51527180",
  1690 => x"2eb33880",
  1691 => x"e1e80852",
  1692 => x"71802e8a",
  1693 => x"38ff1280",
  1694 => x"e1e80cb5",
  1695 => x"9d0480e1",
  1696 => x"e4081080",
  1697 => x"e1e40805",
  1698 => x"70842916",
  1699 => x"51528812",
  1700 => x"08802e89",
  1701 => x"38ff5188",
  1702 => x"12085271",
  1703 => x"2d81f251",
  1704 => x"aca12d80",
  1705 => x"e1840881",
  1706 => x"2a708106",
  1707 => x"51527180",
  1708 => x"2eb43880",
  1709 => x"e1e408ff",
  1710 => x"1180e1e8",
  1711 => x"08565353",
  1712 => x"7372258a",
  1713 => x"38811480",
  1714 => x"e1e80cb5",
  1715 => x"e6047210",
  1716 => x"13708429",
  1717 => x"16515288",
  1718 => x"1208802e",
  1719 => x"8938fe51",
  1720 => x"88120852",
  1721 => x"712d81fd",
  1722 => x"51aca12d",
  1723 => x"80e18408",
  1724 => x"812a7081",
  1725 => x"06515271",
  1726 => x"802eb138",
  1727 => x"80e1e808",
  1728 => x"802e8a38",
  1729 => x"800b80e1",
  1730 => x"e80cb6ac",
  1731 => x"0480e1e4",
  1732 => x"081080e1",
  1733 => x"e4080570",
  1734 => x"84291651",
  1735 => x"52881208",
  1736 => x"802e8938",
  1737 => x"fd518812",
  1738 => x"0852712d",
  1739 => x"81fa51ac",
  1740 => x"a12d80e1",
  1741 => x"8408812a",
  1742 => x"70810651",
  1743 => x"5271802e",
  1744 => x"b13880e1",
  1745 => x"e408ff11",
  1746 => x"545280e1",
  1747 => x"e8087325",
  1748 => x"89387280",
  1749 => x"e1e80cb6",
  1750 => x"f2047110",
  1751 => x"12708429",
  1752 => x"16515288",
  1753 => x"1208802e",
  1754 => x"8938fc51",
  1755 => x"88120852",
  1756 => x"712d80e1",
  1757 => x"e8087053",
  1758 => x"5473802e",
  1759 => x"8a388c15",
  1760 => x"ff155555",
  1761 => x"b6f90482",
  1762 => x"0b80e198",
  1763 => x"0c718f06",
  1764 => x"80e1940c",
  1765 => x"81eb51ac",
  1766 => x"a12d80e1",
  1767 => x"8408812a",
  1768 => x"70810651",
  1769 => x"5271802e",
  1770 => x"ad387408",
  1771 => x"852e0981",
  1772 => x"06a43888",
  1773 => x"1580f52d",
  1774 => x"ff055271",
  1775 => x"881681b7",
  1776 => x"2d71982b",
  1777 => x"52718025",
  1778 => x"8838800b",
  1779 => x"881681b7",
  1780 => x"2d7451af",
  1781 => x"862d81f4",
  1782 => x"51aca12d",
  1783 => x"80e18408",
  1784 => x"812a7081",
  1785 => x"06515271",
  1786 => x"802eb338",
  1787 => x"7408852e",
  1788 => x"098106aa",
  1789 => x"38881580",
  1790 => x"f52d8105",
  1791 => x"52718816",
  1792 => x"81b72d71",
  1793 => x"81ff068b",
  1794 => x"1680f52d",
  1795 => x"54527272",
  1796 => x"27873872",
  1797 => x"881681b7",
  1798 => x"2d7451af",
  1799 => x"862d80da",
  1800 => x"51aca12d",
  1801 => x"80e18408",
  1802 => x"812a7081",
  1803 => x"06515271",
  1804 => x"802e81ad",
  1805 => x"3880e1e0",
  1806 => x"0880e1e8",
  1807 => x"08555373",
  1808 => x"802e8a38",
  1809 => x"8c13ff15",
  1810 => x"5553b8bf",
  1811 => x"04720852",
  1812 => x"71822ea6",
  1813 => x"38718226",
  1814 => x"89387181",
  1815 => x"2eaa38b9",
  1816 => x"e1047183",
  1817 => x"2eb43871",
  1818 => x"842e0981",
  1819 => x"0680f238",
  1820 => x"88130851",
  1821 => x"b0dc2db9",
  1822 => x"e10480e1",
  1823 => x"e8085188",
  1824 => x"13085271",
  1825 => x"2db9e104",
  1826 => x"810b8814",
  1827 => x"082b80df",
  1828 => x"94083280",
  1829 => x"df940cb9",
  1830 => x"b5048813",
  1831 => x"80f52d81",
  1832 => x"058b1480",
  1833 => x"f52d5354",
  1834 => x"71742483",
  1835 => x"38805473",
  1836 => x"881481b7",
  1837 => x"2dafb62d",
  1838 => x"b9e10475",
  1839 => x"08802ea4",
  1840 => x"38750851",
  1841 => x"aca12d80",
  1842 => x"e1840881",
  1843 => x"06527180",
  1844 => x"2e8c3880",
  1845 => x"e1e80851",
  1846 => x"84160852",
  1847 => x"712d8816",
  1848 => x"5675d838",
  1849 => x"8054800b",
  1850 => x"80e1980c",
  1851 => x"738f0680",
  1852 => x"e1940ca0",
  1853 => x"527380e1",
  1854 => x"e8082e09",
  1855 => x"81069938",
  1856 => x"80e1e408",
  1857 => x"ff057432",
  1858 => x"70098105",
  1859 => x"7072079f",
  1860 => x"2a917131",
  1861 => x"51515353",
  1862 => x"71518384",
  1863 => x"2d811454",
  1864 => x"8e7425c2",
  1865 => x"3880df98",
  1866 => x"08527180",
  1867 => x"e1840c02",
  1868 => x"98050d04",
  1869 => x"02f4050d",
  1870 => x"d45281ff",
  1871 => x"720c7108",
  1872 => x"5381ff72",
  1873 => x"0c72882b",
  1874 => x"83fe8006",
  1875 => x"72087081",
  1876 => x"ff065152",
  1877 => x"5381ff72",
  1878 => x"0c727107",
  1879 => x"882b7208",
  1880 => x"7081ff06",
  1881 => x"51525381",
  1882 => x"ff720c72",
  1883 => x"7107882b",
  1884 => x"72087081",
  1885 => x"ff067207",
  1886 => x"80e1840c",
  1887 => x"5253028c",
  1888 => x"050d0402",
  1889 => x"f4050d74",
  1890 => x"767181ff",
  1891 => x"06d40c53",
  1892 => x"5380e1f0",
  1893 => x"08853871",
  1894 => x"892b5271",
  1895 => x"982ad40c",
  1896 => x"71902a70",
  1897 => x"81ff06d4",
  1898 => x"0c517188",
  1899 => x"2a7081ff",
  1900 => x"06d40c51",
  1901 => x"7181ff06",
  1902 => x"d40c7290",
  1903 => x"2a7081ff",
  1904 => x"06d40c51",
  1905 => x"d4087081",
  1906 => x"ff065151",
  1907 => x"82b8bf52",
  1908 => x"7081ff2e",
  1909 => x"09810694",
  1910 => x"3881ff0b",
  1911 => x"d40cd408",
  1912 => x"7081ff06",
  1913 => x"ff145451",
  1914 => x"5171e538",
  1915 => x"7080e184",
  1916 => x"0c028c05",
  1917 => x"0d0402fc",
  1918 => x"050d81c7",
  1919 => x"5181ff0b",
  1920 => x"d40cff11",
  1921 => x"51708025",
  1922 => x"f4380284",
  1923 => x"050d0402",
  1924 => x"f4050d81",
  1925 => x"ff0bd40c",
  1926 => x"93538052",
  1927 => x"87fc80c1",
  1928 => x"51bb832d",
  1929 => x"80e18408",
  1930 => x"8b3881ff",
  1931 => x"0bd40c81",
  1932 => x"53bcbd04",
  1933 => x"bbf62dff",
  1934 => x"135372de",
  1935 => x"387280e1",
  1936 => x"840c028c",
  1937 => x"050d0402",
  1938 => x"ec050d81",
  1939 => x"0b80e1f0",
  1940 => x"0c8454d0",
  1941 => x"08708f2a",
  1942 => x"70810651",
  1943 => x"515372f3",
  1944 => x"3872d00c",
  1945 => x"bbf62d80",
  1946 => x"dad05186",
  1947 => x"a02dd008",
  1948 => x"708f2a70",
  1949 => x"81065151",
  1950 => x"5372f338",
  1951 => x"810bd00c",
  1952 => x"b1538052",
  1953 => x"84d480c0",
  1954 => x"51bb832d",
  1955 => x"80e18408",
  1956 => x"812e9338",
  1957 => x"72822ebf",
  1958 => x"38ff1353",
  1959 => x"72e438ff",
  1960 => x"145473ff",
  1961 => x"ae38bbf6",
  1962 => x"2d83aa52",
  1963 => x"849c80c8",
  1964 => x"51bb832d",
  1965 => x"80e18408",
  1966 => x"812e0981",
  1967 => x"069338ba",
  1968 => x"b42d80e1",
  1969 => x"840883ff",
  1970 => x"ff065372",
  1971 => x"83aa2e9f",
  1972 => x"38bc8f2d",
  1973 => x"bdea0480",
  1974 => x"dadc5186",
  1975 => x"a02d8053",
  1976 => x"bfbf0480",
  1977 => x"daf45186",
  1978 => x"a02d8054",
  1979 => x"bf900481",
  1980 => x"ff0bd40c",
  1981 => x"b154bbf6",
  1982 => x"2d8fcf53",
  1983 => x"805287fc",
  1984 => x"80f751bb",
  1985 => x"832d80e1",
  1986 => x"84085580",
  1987 => x"e1840881",
  1988 => x"2e098106",
  1989 => x"9c3881ff",
  1990 => x"0bd40c82",
  1991 => x"0a52849c",
  1992 => x"80e951bb",
  1993 => x"832d80e1",
  1994 => x"8408802e",
  1995 => x"8d38bbf6",
  1996 => x"2dff1353",
  1997 => x"72c638bf",
  1998 => x"830481ff",
  1999 => x"0bd40c80",
  2000 => x"e1840852",
  2001 => x"87fc80fa",
  2002 => x"51bb832d",
  2003 => x"80e18408",
  2004 => x"b23881ff",
  2005 => x"0bd40cd4",
  2006 => x"085381ff",
  2007 => x"0bd40c81",
  2008 => x"ff0bd40c",
  2009 => x"81ff0bd4",
  2010 => x"0c81ff0b",
  2011 => x"d40c7286",
  2012 => x"2a708106",
  2013 => x"76565153",
  2014 => x"72963880",
  2015 => x"e1840854",
  2016 => x"bf900473",
  2017 => x"822efedb",
  2018 => x"38ff1454",
  2019 => x"73fee738",
  2020 => x"7380e1f0",
  2021 => x"0c738b38",
  2022 => x"815287fc",
  2023 => x"80d051bb",
  2024 => x"832d81ff",
  2025 => x"0bd40cd0",
  2026 => x"08708f2a",
  2027 => x"70810651",
  2028 => x"515372f3",
  2029 => x"3872d00c",
  2030 => x"81ff0bd4",
  2031 => x"0c815372",
  2032 => x"80e1840c",
  2033 => x"0294050d",
  2034 => x"0402e805",
  2035 => x"0d785580",
  2036 => x"5681ff0b",
  2037 => x"d40cd008",
  2038 => x"708f2a70",
  2039 => x"81065151",
  2040 => x"5372f338",
  2041 => x"82810bd0",
  2042 => x"0c81ff0b",
  2043 => x"d40c7752",
  2044 => x"87fc80d1",
  2045 => x"51bb832d",
  2046 => x"80dbc6df",
  2047 => x"5480e184",
  2048 => x"08802e8c",
  2049 => x"3880db94",
  2050 => x"5186a02d",
  2051 => x"80c0e504",
  2052 => x"81ff0bd4",
  2053 => x"0cd40870",
  2054 => x"81ff0651",
  2055 => x"537281fe",
  2056 => x"2e098106",
  2057 => x"9f3880ff",
  2058 => x"53bab42d",
  2059 => x"80e18408",
  2060 => x"75708405",
  2061 => x"570cff13",
  2062 => x"53728025",
  2063 => x"ec388156",
  2064 => x"80c0ca04",
  2065 => x"ff145473",
  2066 => x"c73881ff",
  2067 => x"0bd40c81",
  2068 => x"ff0bd40c",
  2069 => x"d008708f",
  2070 => x"2a708106",
  2071 => x"51515372",
  2072 => x"f33872d0",
  2073 => x"0c7580e1",
  2074 => x"840c0298",
  2075 => x"050d0402",
  2076 => x"e8050d77",
  2077 => x"797b5855",
  2078 => x"55805372",
  2079 => x"7625a538",
  2080 => x"74708105",
  2081 => x"5680f52d",
  2082 => x"74708105",
  2083 => x"5680f52d",
  2084 => x"52527171",
  2085 => x"2e873881",
  2086 => x"5180c1a6",
  2087 => x"04811353",
  2088 => x"80c0fb04",
  2089 => x"80517080",
  2090 => x"e1840c02",
  2091 => x"98050d04",
  2092 => x"02ec050d",
  2093 => x"76557480",
  2094 => x"2e80c438",
  2095 => x"9a1580e0",
  2096 => x"2d5180d1",
  2097 => x"8e2d80e1",
  2098 => x"840880e1",
  2099 => x"840880e8",
  2100 => x"a40c80e1",
  2101 => x"84085454",
  2102 => x"80e88008",
  2103 => x"802e9b38",
  2104 => x"941580e0",
  2105 => x"2d5180d1",
  2106 => x"8e2d80e1",
  2107 => x"8408902b",
  2108 => x"83fff00a",
  2109 => x"06707507",
  2110 => x"51537280",
  2111 => x"e8a40c80",
  2112 => x"e8a40853",
  2113 => x"72802e9e",
  2114 => x"3880e7f8",
  2115 => x"08fe1471",
  2116 => x"2980e88c",
  2117 => x"080580e8",
  2118 => x"a80c7084",
  2119 => x"2b80e884",
  2120 => x"0c5480c2",
  2121 => x"d50480e8",
  2122 => x"900880e8",
  2123 => x"a40c80e8",
  2124 => x"940880e8",
  2125 => x"a80c80e8",
  2126 => x"8008802e",
  2127 => x"8c3880e7",
  2128 => x"f808842b",
  2129 => x"5380c2d0",
  2130 => x"0480e898",
  2131 => x"08842b53",
  2132 => x"7280e884",
  2133 => x"0c029405",
  2134 => x"0d0402d8",
  2135 => x"050d800b",
  2136 => x"80e8800c",
  2137 => x"8454bcc7",
  2138 => x"2d80e184",
  2139 => x"08802e98",
  2140 => x"3880e1f4",
  2141 => x"528051bf",
  2142 => x"c92d80e1",
  2143 => x"8408802e",
  2144 => x"8738fe54",
  2145 => x"80c39004",
  2146 => x"ff145473",
  2147 => x"8024d738",
  2148 => x"738e3880",
  2149 => x"dba45186",
  2150 => x"a02d7355",
  2151 => x"80c8f304",
  2152 => x"8056810b",
  2153 => x"80e8ac0c",
  2154 => x"885380db",
  2155 => x"b85280e2",
  2156 => x"aa5180c0",
  2157 => x"ef2d80e1",
  2158 => x"8408762e",
  2159 => x"09810689",
  2160 => x"3880e184",
  2161 => x"0880e8ac",
  2162 => x"0c885380",
  2163 => x"dbc45280",
  2164 => x"e2c65180",
  2165 => x"c0ef2d80",
  2166 => x"e1840889",
  2167 => x"3880e184",
  2168 => x"0880e8ac",
  2169 => x"0c80e8ac",
  2170 => x"08802e81",
  2171 => x"843880e5",
  2172 => x"ba0b80f5",
  2173 => x"2d80e5bb",
  2174 => x"0b80f52d",
  2175 => x"71982b71",
  2176 => x"902b0780",
  2177 => x"e5bc0b80",
  2178 => x"f52d7088",
  2179 => x"2b720780",
  2180 => x"e5bd0b80",
  2181 => x"f52d7107",
  2182 => x"80e5f20b",
  2183 => x"80f52d80",
  2184 => x"e5f30b80",
  2185 => x"f52d7188",
  2186 => x"2b07535f",
  2187 => x"54525a56",
  2188 => x"57557381",
  2189 => x"abaa2e09",
  2190 => x"81069038",
  2191 => x"755180d0",
  2192 => x"dd2d80e1",
  2193 => x"84085680",
  2194 => x"c4da0473",
  2195 => x"82d4d52e",
  2196 => x"893880db",
  2197 => x"d05180c5",
  2198 => x"a90480e1",
  2199 => x"f4527551",
  2200 => x"bfc92d80",
  2201 => x"e1840855",
  2202 => x"80e18408",
  2203 => x"802e8483",
  2204 => x"38885380",
  2205 => x"dbc45280",
  2206 => x"e2c65180",
  2207 => x"c0ef2d80",
  2208 => x"e184088b",
  2209 => x"38810b80",
  2210 => x"e8800c80",
  2211 => x"c5b00488",
  2212 => x"5380dbb8",
  2213 => x"5280e2aa",
  2214 => x"5180c0ef",
  2215 => x"2d80e184",
  2216 => x"08802e8c",
  2217 => x"3880dbe4",
  2218 => x"5186a02d",
  2219 => x"80c68f04",
  2220 => x"80e5f20b",
  2221 => x"80f52d54",
  2222 => x"7380d52e",
  2223 => x"09810680",
  2224 => x"ce3880e5",
  2225 => x"f30b80f5",
  2226 => x"2d547381",
  2227 => x"aa2e0981",
  2228 => x"06bd3880",
  2229 => x"0b80e1f4",
  2230 => x"0b80f52d",
  2231 => x"56547481",
  2232 => x"e92e8338",
  2233 => x"81547481",
  2234 => x"eb2e8c38",
  2235 => x"80557375",
  2236 => x"2e098106",
  2237 => x"82fd3880",
  2238 => x"e1ff0b80",
  2239 => x"f52d5574",
  2240 => x"8e3880e2",
  2241 => x"800b80f5",
  2242 => x"2d547382",
  2243 => x"2e873880",
  2244 => x"5580c8f3",
  2245 => x"0480e281",
  2246 => x"0b80f52d",
  2247 => x"7080e7f8",
  2248 => x"0cff0580",
  2249 => x"e7fc0c80",
  2250 => x"e2820b80",
  2251 => x"f52d80e2",
  2252 => x"830b80f5",
  2253 => x"2d587605",
  2254 => x"77828029",
  2255 => x"057080e8",
  2256 => x"880c80e2",
  2257 => x"840b80f5",
  2258 => x"2d7080e8",
  2259 => x"9c0c80e8",
  2260 => x"80085957",
  2261 => x"5876802e",
  2262 => x"81b93888",
  2263 => x"5380dbc4",
  2264 => x"5280e2c6",
  2265 => x"5180c0ef",
  2266 => x"2d80e184",
  2267 => x"08828438",
  2268 => x"80e7f808",
  2269 => x"70842b80",
  2270 => x"e8840c70",
  2271 => x"80e8980c",
  2272 => x"80e2990b",
  2273 => x"80f52d80",
  2274 => x"e2980b80",
  2275 => x"f52d7182",
  2276 => x"80290580",
  2277 => x"e29a0b80",
  2278 => x"f52d7084",
  2279 => x"80802912",
  2280 => x"80e29b0b",
  2281 => x"80f52d70",
  2282 => x"81800a29",
  2283 => x"127080e8",
  2284 => x"a00c80e8",
  2285 => x"9c087129",
  2286 => x"80e88808",
  2287 => x"057080e8",
  2288 => x"8c0c80e2",
  2289 => x"a10b80f5",
  2290 => x"2d80e2a0",
  2291 => x"0b80f52d",
  2292 => x"71828029",
  2293 => x"0580e2a2",
  2294 => x"0b80f52d",
  2295 => x"70848080",
  2296 => x"291280e2",
  2297 => x"a30b80f5",
  2298 => x"2d70982b",
  2299 => x"81f00a06",
  2300 => x"72057080",
  2301 => x"e8900cfe",
  2302 => x"117e2977",
  2303 => x"0580e894",
  2304 => x"0c525952",
  2305 => x"43545e51",
  2306 => x"5259525d",
  2307 => x"57595780",
  2308 => x"c8eb0480",
  2309 => x"e2860b80",
  2310 => x"f52d80e2",
  2311 => x"850b80f5",
  2312 => x"2d718280",
  2313 => x"29057080",
  2314 => x"e8840c70",
  2315 => x"a02983ff",
  2316 => x"0570892a",
  2317 => x"7080e898",
  2318 => x"0c80e28b",
  2319 => x"0b80f52d",
  2320 => x"80e28a0b",
  2321 => x"80f52d71",
  2322 => x"82802905",
  2323 => x"7080e8a0",
  2324 => x"0c7b7129",
  2325 => x"1e7080e8",
  2326 => x"940c7d80",
  2327 => x"e8900c73",
  2328 => x"0580e88c",
  2329 => x"0c555e51",
  2330 => x"51555580",
  2331 => x"5180c1b0",
  2332 => x"2d815574",
  2333 => x"80e1840c",
  2334 => x"02a8050d",
  2335 => x"0402ec05",
  2336 => x"0d767087",
  2337 => x"2c7180ff",
  2338 => x"06555654",
  2339 => x"80e88008",
  2340 => x"8a387388",
  2341 => x"2c7481ff",
  2342 => x"06545580",
  2343 => x"e1f45280",
  2344 => x"e8880815",
  2345 => x"51bfc92d",
  2346 => x"80e18408",
  2347 => x"5480e184",
  2348 => x"08802ebb",
  2349 => x"3880e880",
  2350 => x"08802e9c",
  2351 => x"38728429",
  2352 => x"80e1f405",
  2353 => x"70085253",
  2354 => x"80d0dd2d",
  2355 => x"80e18408",
  2356 => x"f00a0653",
  2357 => x"80c9ed04",
  2358 => x"721080e1",
  2359 => x"f4057080",
  2360 => x"e02d5253",
  2361 => x"80d18e2d",
  2362 => x"80e18408",
  2363 => x"53725473",
  2364 => x"80e1840c",
  2365 => x"0294050d",
  2366 => x"0402e005",
  2367 => x"0d797b59",
  2368 => x"54805577",
  2369 => x"752e8438",
  2370 => x"74780c73",
  2371 => x"842c80e8",
  2372 => x"a8080574",
  2373 => x"8f065457",
  2374 => x"72818038",
  2375 => x"80e88008",
  2376 => x"802e80ee",
  2377 => x"3880e8a4",
  2378 => x"085680e8",
  2379 => x"84087426",
  2380 => x"80d83875",
  2381 => x"5180c8fd",
  2382 => x"2d80e184",
  2383 => x"0880e184",
  2384 => x"0880ffff",
  2385 => x"fff80654",
  2386 => x"567280ff",
  2387 => x"fffff82e",
  2388 => x"83813880",
  2389 => x"e8840874",
  2390 => x"71318117",
  2391 => x"57555373",
  2392 => x"7327d038",
  2393 => x"74802ea2",
  2394 => x"3880e184",
  2395 => x"08fe0580",
  2396 => x"e7f80829",
  2397 => x"80e88c08",
  2398 => x"0574842c",
  2399 => x"0580e184",
  2400 => x"0880df9c",
  2401 => x"0c5780cb",
  2402 => x"920480e8",
  2403 => x"a40880df",
  2404 => x"9c0c80e1",
  2405 => x"f4527651",
  2406 => x"bfc92d73",
  2407 => x"852b83e0",
  2408 => x"0680e1f4",
  2409 => x"05558075",
  2410 => x"80f52d54",
  2411 => x"5672762e",
  2412 => x"09810683",
  2413 => x"38815677",
  2414 => x"802e8f38",
  2415 => x"81707706",
  2416 => x"54547280",
  2417 => x"2e843873",
  2418 => x"780c8075",
  2419 => x"80f52d55",
  2420 => x"5373732e",
  2421 => x"83388153",
  2422 => x"7381e52e",
  2423 => x"81f53881",
  2424 => x"70740654",
  2425 => x"5872802e",
  2426 => x"81e9388b",
  2427 => x"1580f52d",
  2428 => x"70832a79",
  2429 => x"06585676",
  2430 => x"9c3880df",
  2431 => x"a0085372",
  2432 => x"89387280",
  2433 => x"e5f40b81",
  2434 => x"b72d7680",
  2435 => x"dfa00c74",
  2436 => x"5380cdd5",
  2437 => x"04758f2e",
  2438 => x"09810681",
  2439 => x"b638739f",
  2440 => x"068d2980",
  2441 => x"e5e71151",
  2442 => x"53811580",
  2443 => x"f52d7370",
  2444 => x"81055581",
  2445 => x"b72d8315",
  2446 => x"80f52d73",
  2447 => x"70810555",
  2448 => x"81b72d85",
  2449 => x"1580f52d",
  2450 => x"73708105",
  2451 => x"5581b72d",
  2452 => x"871580f5",
  2453 => x"2d737081",
  2454 => x"055581b7",
  2455 => x"2d891580",
  2456 => x"f52d7370",
  2457 => x"81055581",
  2458 => x"b72d8e15",
  2459 => x"80f52d73",
  2460 => x"70810555",
  2461 => x"81b72d90",
  2462 => x"1580f52d",
  2463 => x"73708105",
  2464 => x"5581b72d",
  2465 => x"921580f5",
  2466 => x"2d737081",
  2467 => x"055581b7",
  2468 => x"2d941580",
  2469 => x"f52d7370",
  2470 => x"81055581",
  2471 => x"b72d9615",
  2472 => x"80f52d73",
  2473 => x"70810555",
  2474 => x"81b72d98",
  2475 => x"1580f52d",
  2476 => x"73708105",
  2477 => x"5581b72d",
  2478 => x"9c1580f5",
  2479 => x"2d737081",
  2480 => x"055581b7",
  2481 => x"2d9e1580",
  2482 => x"f52d7381",
  2483 => x"b72d7780",
  2484 => x"dfa00c80",
  2485 => x"537280e1",
  2486 => x"840c02a0",
  2487 => x"050d0402",
  2488 => x"cc050d7e",
  2489 => x"605e5a80",
  2490 => x"0b80e8a4",
  2491 => x"0880e8a8",
  2492 => x"08595c56",
  2493 => x"805880e8",
  2494 => x"8408782e",
  2495 => x"81bd3877",
  2496 => x"8f06a017",
  2497 => x"57547391",
  2498 => x"3880e1f4",
  2499 => x"52765181",
  2500 => x"1757bfc9",
  2501 => x"2d80e1f4",
  2502 => x"56807680",
  2503 => x"f52d5654",
  2504 => x"74742e83",
  2505 => x"38815474",
  2506 => x"81e52e81",
  2507 => x"82388170",
  2508 => x"7506555c",
  2509 => x"73802e80",
  2510 => x"f6388b16",
  2511 => x"80f52d98",
  2512 => x"06597880",
  2513 => x"ea388b53",
  2514 => x"7c527551",
  2515 => x"80c0ef2d",
  2516 => x"80e18408",
  2517 => x"80d9389c",
  2518 => x"16085180",
  2519 => x"d0dd2d80",
  2520 => x"e1840884",
  2521 => x"1b0c9a16",
  2522 => x"80e02d51",
  2523 => x"80d18e2d",
  2524 => x"80e18408",
  2525 => x"80e18408",
  2526 => x"881c0c80",
  2527 => x"e1840855",
  2528 => x"5580e880",
  2529 => x"08802e9a",
  2530 => x"38941680",
  2531 => x"e02d5180",
  2532 => x"d18e2d80",
  2533 => x"e1840890",
  2534 => x"2b83fff0",
  2535 => x"0a067016",
  2536 => x"51547388",
  2537 => x"1b0c787a",
  2538 => x"0c7b5480",
  2539 => x"cff90481",
  2540 => x"185880e8",
  2541 => x"84087826",
  2542 => x"fec53880",
  2543 => x"e8800880",
  2544 => x"2eb5387a",
  2545 => x"5180c8fd",
  2546 => x"2d80e184",
  2547 => x"0880e184",
  2548 => x"0880ffff",
  2549 => x"fff80655",
  2550 => x"5b7380ff",
  2551 => x"fffff82e",
  2552 => x"963880e1",
  2553 => x"8408fe05",
  2554 => x"80e7f808",
  2555 => x"2980e88c",
  2556 => x"08055780",
  2557 => x"cdf40480",
  2558 => x"547380e1",
  2559 => x"840c02b4",
  2560 => x"050d0402",
  2561 => x"f4050d74",
  2562 => x"70088105",
  2563 => x"710c7008",
  2564 => x"80e7fc08",
  2565 => x"06535371",
  2566 => x"90388813",
  2567 => x"085180c8",
  2568 => x"fd2d80e1",
  2569 => x"84088814",
  2570 => x"0c810b80",
  2571 => x"e1840c02",
  2572 => x"8c050d04",
  2573 => x"02f0050d",
  2574 => x"75881108",
  2575 => x"fe0580e7",
  2576 => x"f8082980",
  2577 => x"e88c0811",
  2578 => x"720880e7",
  2579 => x"fc080605",
  2580 => x"79555354",
  2581 => x"54bfc92d",
  2582 => x"0290050d",
  2583 => x"0402f405",
  2584 => x"0d747088",
  2585 => x"2a83fe80",
  2586 => x"06707298",
  2587 => x"2a077288",
  2588 => x"2b87fc80",
  2589 => x"80067398",
  2590 => x"2b81f00a",
  2591 => x"06717307",
  2592 => x"0780e184",
  2593 => x"0c565153",
  2594 => x"51028c05",
  2595 => x"0d0402f8",
  2596 => x"050d028e",
  2597 => x"0580f52d",
  2598 => x"74882b07",
  2599 => x"7083ffff",
  2600 => x"0680e184",
  2601 => x"0c510288",
  2602 => x"050d0402",
  2603 => x"f4050d74",
  2604 => x"76785354",
  2605 => x"52807125",
  2606 => x"97387270",
  2607 => x"81055480",
  2608 => x"f52d7270",
  2609 => x"81055481",
  2610 => x"b72dff11",
  2611 => x"5170eb38",
  2612 => x"807281b7",
  2613 => x"2d028c05",
  2614 => x"0d0402e0",
  2615 => x"050d7957",
  2616 => x"80705970",
  2617 => x"575580d2",
  2618 => x"910402a0",
  2619 => x"05fc0552",
  2620 => x"755180c9",
  2621 => x"f92d80e1",
  2622 => x"840880e1",
  2623 => x"84080981",
  2624 => x"057080e1",
  2625 => x"8408079f",
  2626 => x"2a770581",
  2627 => x"19595754",
  2628 => x"54767525",
  2629 => x"53778438",
  2630 => x"72d03873",
  2631 => x"80e1840c",
  2632 => x"02a0050d",
  2633 => x"0402f005",
  2634 => x"0d80e180",
  2635 => x"08165180",
  2636 => x"d1da2d80",
  2637 => x"e1840880",
  2638 => x"2ea0388b",
  2639 => x"5380e184",
  2640 => x"085280e5",
  2641 => x"f45180d1",
  2642 => x"ab2d80e8",
  2643 => x"b0085473",
  2644 => x"802e8738",
  2645 => x"80e5f451",
  2646 => x"732d0290",
  2647 => x"050d0402",
  2648 => x"f4050d74",
  2649 => x"76708c2c",
  2650 => x"708f0680",
  2651 => x"dc940805",
  2652 => x"51535353",
  2653 => x"7080f52d",
  2654 => x"7381b72d",
  2655 => x"71882c70",
  2656 => x"8f0680dc",
  2657 => x"94080551",
  2658 => x"517080f5",
  2659 => x"2d811481",
  2660 => x"b72d7184",
  2661 => x"2c708f06",
  2662 => x"80dc9408",
  2663 => x"05515170",
  2664 => x"80f52d82",
  2665 => x"1481b72d",
  2666 => x"718f0680",
  2667 => x"dc940805",
  2668 => x"527180f5",
  2669 => x"2d831481",
  2670 => x"b72d028c",
  2671 => x"050d0402",
  2672 => x"d8050d80",
  2673 => x"5a807056",
  2674 => x"5980d3ef",
  2675 => x"0402a805",
  2676 => x"fc055278",
  2677 => x"5180c9f9",
  2678 => x"2d80e184",
  2679 => x"08098105",
  2680 => x"7080e184",
  2681 => x"08079f2a",
  2682 => x"7605811b",
  2683 => x"5b565480",
  2684 => x"e1800875",
  2685 => x"24547984",
  2686 => x"3873d238",
  2687 => x"80705b55",
  2688 => x"02a805fc",
  2689 => x"05527851",
  2690 => x"80c9f92d",
  2691 => x"80e18408",
  2692 => x"802e81b4",
  2693 => x"3880e184",
  2694 => x"088b0580",
  2695 => x"f52d7084",
  2696 => x"2a708106",
  2697 => x"77107884",
  2698 => x"2b80e5f4",
  2699 => x"0b80f52d",
  2700 => x"5c5c5351",
  2701 => x"55567380",
  2702 => x"2e80ce38",
  2703 => x"7416822b",
  2704 => x"80d7de0b",
  2705 => x"80dfac12",
  2706 => x"0c547775",
  2707 => x"311080e8",
  2708 => x"b4115556",
  2709 => x"90747081",
  2710 => x"055681b7",
  2711 => x"2da07481",
  2712 => x"b72d7681",
  2713 => x"ff068116",
  2714 => x"58547380",
  2715 => x"2e8b389c",
  2716 => x"5380e5f4",
  2717 => x"5280d580",
  2718 => x"048b5380",
  2719 => x"e1840852",
  2720 => x"80e8b616",
  2721 => x"5180d5be",
  2722 => x"04741682",
  2723 => x"2b80d2a5",
  2724 => x"0b80dfac",
  2725 => x"120c5476",
  2726 => x"81ff0681",
  2727 => x"16585473",
  2728 => x"802e8b38",
  2729 => x"9c5380e5",
  2730 => x"f45280d5",
  2731 => x"b5048b53",
  2732 => x"80e18408",
  2733 => x"52777531",
  2734 => x"1080e8b4",
  2735 => x"05517655",
  2736 => x"80d1ab2d",
  2737 => x"80d5dd04",
  2738 => x"74902975",
  2739 => x"31701080",
  2740 => x"e8b40551",
  2741 => x"5480e184",
  2742 => x"087481b7",
  2743 => x"2d811959",
  2744 => x"748b24a6",
  2745 => x"3879802e",
  2746 => x"fe963874",
  2747 => x"90297531",
  2748 => x"701080e8",
  2749 => x"b4058c77",
  2750 => x"31575154",
  2751 => x"807481b7",
  2752 => x"2d9e14ff",
  2753 => x"16565474",
  2754 => x"f33880db",
  2755 => x"f05280e0",
  2756 => x"d851a290",
  2757 => x"2d80e180",
  2758 => x"085280e0",
  2759 => x"dd5180d2",
  2760 => x"df2d80e8",
  2761 => x"84085280",
  2762 => x"e0e25180",
  2763 => x"d2df2d78",
  2764 => x"5280e0e7",
  2765 => x"5180d2df",
  2766 => x"2d80df9c",
  2767 => x"0b80e02d",
  2768 => x"5280e0ec",
  2769 => x"5180d2df",
  2770 => x"2d80df9e",
  2771 => x"0b80e02d",
  2772 => x"5280e0f0",
  2773 => x"5180d2df",
  2774 => x"2d7880e1",
  2775 => x"840c02a8",
  2776 => x"050d0402",
  2777 => x"fc050d72",
  2778 => x"5170fd2e",
  2779 => x"b23870fd",
  2780 => x"248b3870",
  2781 => x"fc2e80d0",
  2782 => x"3880d7d2",
  2783 => x"0470fe2e",
  2784 => x"b93870ff",
  2785 => x"2e098106",
  2786 => x"80c83880",
  2787 => x"e1800851",
  2788 => x"70802ebe",
  2789 => x"38ff1180",
  2790 => x"e1800c80",
  2791 => x"d7d20480",
  2792 => x"e18008f4",
  2793 => x"057080e1",
  2794 => x"800c5170",
  2795 => x"8025a338",
  2796 => x"800b80e1",
  2797 => x"800c80d7",
  2798 => x"d20480e1",
  2799 => x"80088105",
  2800 => x"80e1800c",
  2801 => x"80d7d204",
  2802 => x"80e18008",
  2803 => x"8c0580e1",
  2804 => x"800c80d3",
  2805 => x"bf2dafb6",
  2806 => x"2d028405",
  2807 => x"0d0402fc",
  2808 => x"050d80e1",
  2809 => x"80081351",
  2810 => x"80d1da2d",
  2811 => x"80e18408",
  2812 => x"802e8a38",
  2813 => x"80e18408",
  2814 => x"5180c1b0",
  2815 => x"2d800b80",
  2816 => x"e1800c80",
  2817 => x"d3bf2daf",
  2818 => x"b62d0284",
  2819 => x"050d0402",
  2820 => x"fc050d80",
  2821 => x"0b80e180",
  2822 => x"0c80d3bf",
  2823 => x"2daeb22d",
  2824 => x"80e18408",
  2825 => x"80e0c80c",
  2826 => x"80dfa451",
  2827 => x"b0dc2d02",
  2828 => x"84050d04",
  2829 => x"7180e8b0",
  2830 => x"0c040000",
  2831 => x"00ffffff",
  2832 => x"ff00ffff",
  2833 => x"ffff00ff",
  2834 => x"ffffff00",
  2835 => x"30313233",
  2836 => x"34353637",
  2837 => x"38394142",
  2838 => x"43444546",
  2839 => x"00000000",
  2840 => x"52657365",
  2841 => x"74000000",
  2842 => x"5363616e",
  2843 => x"6c696e65",
  2844 => x"73000000",
  2845 => x"50414c20",
  2846 => x"2f204e54",
  2847 => x"53430000",
  2848 => x"436f6c6f",
  2849 => x"72000000",
  2850 => x"44696666",
  2851 => x"6963756c",
  2852 => x"74792041",
  2853 => x"00000000",
  2854 => x"44696666",
  2855 => x"6963756c",
  2856 => x"74792042",
  2857 => x"00000000",
  2858 => x"2a537570",
  2859 => x"65726368",
  2860 => x"69702069",
  2861 => x"6e206361",
  2862 => x"72747269",
  2863 => x"64676500",
  2864 => x"2a42616e",
  2865 => x"6b204530",
  2866 => x"00000000",
  2867 => x"2a42616e",
  2868 => x"6b204537",
  2869 => x"00000000",
  2870 => x"53656c65",
  2871 => x"63740000",
  2872 => x"53746172",
  2873 => x"74000000",
  2874 => x"4c6f6164",
  2875 => x"20524f4d",
  2876 => x"20100000",
  2877 => x"45786974",
  2878 => x"00000000",
  2879 => x"524f4d20",
  2880 => x"6c6f6164",
  2881 => x"696e6720",
  2882 => x"6661696c",
  2883 => x"65640000",
  2884 => x"4f4b0000",
  2885 => x"496e6974",
  2886 => x"69616c69",
  2887 => x"7a696e67",
  2888 => x"20534420",
  2889 => x"63617264",
  2890 => x"0a000000",
  2891 => x"446f6e65",
  2892 => x"20696e69",
  2893 => x"7469616c",
  2894 => x"697a6174",
  2895 => x"696f6e0a",
  2896 => x"00000000",
  2897 => x"16200000",
  2898 => x"14200000",
  2899 => x"15200000",
  2900 => x"53442069",
  2901 => x"6e69742e",
  2902 => x"2e2e0a00",
  2903 => x"53442063",
  2904 => x"61726420",
  2905 => x"72657365",
  2906 => x"74206661",
  2907 => x"696c6564",
  2908 => x"210a0000",
  2909 => x"53444843",
  2910 => x"20657272",
  2911 => x"6f72210a",
  2912 => x"00000000",
  2913 => x"57726974",
  2914 => x"65206661",
  2915 => x"696c6564",
  2916 => x"0a000000",
  2917 => x"52656164",
  2918 => x"20666169",
  2919 => x"6c65640a",
  2920 => x"00000000",
  2921 => x"43617264",
  2922 => x"20696e69",
  2923 => x"74206661",
  2924 => x"696c6564",
  2925 => x"0a000000",
  2926 => x"46415431",
  2927 => x"36202020",
  2928 => x"00000000",
  2929 => x"46415433",
  2930 => x"32202020",
  2931 => x"00000000",
  2932 => x"4e6f2070",
  2933 => x"61727469",
  2934 => x"74696f6e",
  2935 => x"20736967",
  2936 => x"0a000000",
  2937 => x"42616420",
  2938 => x"70617274",
  2939 => x"0a000000",
  2940 => x"4261636b",
  2941 => x"20787878",
  2942 => x"78207979",
  2943 => x"7979207a",
  2944 => x"7a7a7a20",
  2945 => x"6b6b6b6b",
  2946 => x"6b6b6b6b",
  2947 => x"00000000",
  2948 => x"00000002",
  2949 => x"00002c4c",
  2950 => x"00000002",
  2951 => x"00002c60",
  2952 => x"0000035a",
  2953 => x"00000001",
  2954 => x"00002c68",
  2955 => x"00000000",
  2956 => x"00000001",
  2957 => x"00002c74",
  2958 => x"00000001",
  2959 => x"00000001",
  2960 => x"00002c80",
  2961 => x"00000002",
  2962 => x"00000001",
  2963 => x"00002c88",
  2964 => x"00000003",
  2965 => x"00000001",
  2966 => x"00002c98",
  2967 => x"00000004",
  2968 => x"00000001",
  2969 => x"00002ca8",
  2970 => x"00000005",
  2971 => x"00000001",
  2972 => x"00002cc0",
  2973 => x"00000008",
  2974 => x"00000001",
  2975 => x"00002ccc",
  2976 => x"00000009",
  2977 => x"00000002",
  2978 => x"00002cd8",
  2979 => x"0000036e",
  2980 => x"00000002",
  2981 => x"00002ce0",
  2982 => x"00000a3f",
  2983 => x"00000002",
  2984 => x"00002ce8",
  2985 => x"00002c0f",
  2986 => x"00000002",
  2987 => x"00002cf4",
  2988 => x"0000174f",
  2989 => x"00000000",
  2990 => x"00000000",
  2991 => x"00000000",
  2992 => x"00000004",
  2993 => x"00002cfc",
  2994 => x"00002ec0",
  2995 => x"00000004",
  2996 => x"00002d10",
  2997 => x"00002e18",
  2998 => x"00000000",
  2999 => x"00000000",
  3000 => x"00000000",
  3001 => x"00000000",
  3002 => x"00000000",
  3003 => x"00000000",
  3004 => x"00000000",
  3005 => x"00000000",
  3006 => x"00000000",
  3007 => x"00000000",
  3008 => x"00000000",
  3009 => x"00000000",
  3010 => x"00000000",
  3011 => x"00000000",
  3012 => x"00000000",
  3013 => x"00000000",
  3014 => x"00000000",
  3015 => x"00000000",
  3016 => x"00000000",
  3017 => x"761c1c1c",
  3018 => x"1c1c051c",
  3019 => x"1c1c1c1c",
  3020 => x"f2f5fafd",
  3021 => x"5a000000",
  3022 => x"00000000",
  3023 => x"00000000",
  3024 => x"00000000",
  3025 => x"00000000",
  3026 => x"00000000",
  3027 => x"00000000",
  3028 => x"00000000",
  3029 => x"00000000",
  3030 => x"00000000",
  3031 => x"00000000",
  3032 => x"00000000",
  3033 => x"00000000",
  3034 => x"00000000",
  3035 => x"00000000",
  3036 => x"00000000",
  3037 => x"00000000",
  3038 => x"00000000",
  3039 => x"00000000",
  3040 => x"0001ffff",
  3041 => x"0001ffff",
  3042 => x"0001ffff",
  3043 => x"00000000",
  3044 => x"00000000",
  3045 => x"00000004",
  3046 => x"00000000",
  3047 => x"00000000",
  3048 => x"00000000",
  3049 => x"00000002",
  3050 => x"00003434",
  3051 => x"00002925",
  3052 => x"00000002",
  3053 => x"00003452",
  3054 => x"00002925",
  3055 => x"00000002",
  3056 => x"00003470",
  3057 => x"00002925",
  3058 => x"00000002",
  3059 => x"0000348e",
  3060 => x"00002925",
  3061 => x"00000002",
  3062 => x"000034ac",
  3063 => x"00002925",
  3064 => x"00000002",
  3065 => x"000034ca",
  3066 => x"00002925",
  3067 => x"00000002",
  3068 => x"000034e8",
  3069 => x"00002925",
  3070 => x"00000002",
  3071 => x"00003506",
  3072 => x"00002925",
  3073 => x"00000002",
  3074 => x"00003524",
  3075 => x"00002925",
  3076 => x"00000002",
  3077 => x"00003542",
  3078 => x"00002925",
  3079 => x"00000002",
  3080 => x"00003560",
  3081 => x"00002925",
  3082 => x"00000002",
  3083 => x"0000357e",
  3084 => x"00002925",
  3085 => x"00000002",
  3086 => x"0000359c",
  3087 => x"00002925",
  3088 => x"00000004",
  3089 => x"00003058",
  3090 => x"00000000",
  3091 => x"00000000",
  3092 => x"00000000",
  3093 => x"00002b63",
  3094 => x"4261636b",
  3095 => x"00000000",
  3096 => x"00000000",
  3097 => x"00000000",
  3098 => x"00000000",
  3099 => x"00000000",
  3100 => x"00000000",
  3101 => x"00000000",
  3102 => x"00000000",
  3103 => x"00000000",
  3104 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

