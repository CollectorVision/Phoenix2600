-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80db",
     9 => x"d0080b0b",
    10 => x"80dbd408",
    11 => x"0b0b80db",
    12 => x"d8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"dbd80c0b",
    16 => x"0b80dbd4",
    17 => x"0c0b0b80",
    18 => x"dbd00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d498",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80dbd070",
    57 => x"80e79027",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a794",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80db",
    65 => x"e00c9f0b",
    66 => x"80dbe40c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"dbe408ff",
    70 => x"0580dbe4",
    71 => x"0c80dbe4",
    72 => x"088025e8",
    73 => x"3880dbe0",
    74 => x"08ff0580",
    75 => x"dbe00c80",
    76 => x"dbe00880",
    77 => x"25d03880",
    78 => x"0b80dbe4",
    79 => x"0c800b80",
    80 => x"dbe00c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80dbe008",
   100 => x"25913882",
   101 => x"c82d80db",
   102 => x"e008ff05",
   103 => x"80dbe00c",
   104 => x"838a0480",
   105 => x"dbe00880",
   106 => x"dbe40853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80dbe008",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"dbe40881",
   116 => x"0580dbe4",
   117 => x"0c80dbe4",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80dbe4",
   121 => x"0c80dbe0",
   122 => x"08810580",
   123 => x"dbe00c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480db",
   128 => x"e4088105",
   129 => x"80dbe40c",
   130 => x"80dbe408",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80dbe4",
   134 => x"0c80dbe0",
   135 => x"08810580",
   136 => x"dbe00c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"dbe80cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"dbe80c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280db",
   177 => x"e8088407",
   178 => x"80dbe80c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80d7",
   183 => x"d00c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80dbe8",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80db",
   208 => x"d00c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02f8050d",
  1093 => x"80da8c08",
  1094 => x"862a7083",
  1095 => x"068207e0",
  1096 => x"0c528051",
  1097 => x"86da2d86",
  1098 => x"c72d0288",
  1099 => x"050d0402",
  1100 => x"f8050d02",
  1101 => x"8f0580f5",
  1102 => x"2d80d7d8",
  1103 => x"08525270",
  1104 => x"80dcfd27",
  1105 => x"9a387171",
  1106 => x"81b72d80",
  1107 => x"d7d80881",
  1108 => x"0580d7d8",
  1109 => x"0c80d7d8",
  1110 => x"08518071",
  1111 => x"81b72d02",
  1112 => x"88050d04",
  1113 => x"02f4050d",
  1114 => x"7470842a",
  1115 => x"708f0680",
  1116 => x"d7d40805",
  1117 => x"7080f52d",
  1118 => x"54515353",
  1119 => x"a2af2d72",
  1120 => x"8f0680d7",
  1121 => x"d4080570",
  1122 => x"80f52d52",
  1123 => x"53a2af2d",
  1124 => x"028c050d",
  1125 => x"0402f405",
  1126 => x"0d747654",
  1127 => x"52727081",
  1128 => x"055480f5",
  1129 => x"2d517072",
  1130 => x"70810554",
  1131 => x"81b72d70",
  1132 => x"ec387072",
  1133 => x"81b72d02",
  1134 => x"8c050d04",
  1135 => x"02c0050d",
  1136 => x"6140800b",
  1137 => x"80da8c08",
  1138 => x"81800671",
  1139 => x"725a4040",
  1140 => x"58810bec",
  1141 => x"0c840bec",
  1142 => x"0c7f5280",
  1143 => x"dbec5180",
  1144 => x"cae72d80",
  1145 => x"dbd00878",
  1146 => x"2e828138",
  1147 => x"80dbf008",
  1148 => x"78ff1257",
  1149 => x"5e567478",
  1150 => x"2e8b3881",
  1151 => x"1d75812a",
  1152 => x"565d74f7",
  1153 => x"38f71d5d",
  1154 => x"81588076",
  1155 => x"2581dd38",
  1156 => x"7c527451",
  1157 => x"84a82d80",
  1158 => x"ddc85280",
  1159 => x"dbec5180",
  1160 => x"cdbb2d80",
  1161 => x"dbd00880",
  1162 => x"2e81a738",
  1163 => x"80ddc85c",
  1164 => x"83ff597e",
  1165 => x"9c387b70",
  1166 => x"81055d80",
  1167 => x"f52d7781",
  1168 => x"1959e40c",
  1169 => x"e80cff19",
  1170 => x"59788025",
  1171 => x"e938a5da",
  1172 => x"047b7081",
  1173 => x"055d80f5",
  1174 => x"2d778119",
  1175 => x"59e40cf4",
  1176 => x"80087072",
  1177 => x"32700981",
  1178 => x"05707207",
  1179 => x"9f2a5156",
  1180 => x"565c5a7d",
  1181 => x"80d03881",
  1182 => x"70740654",
  1183 => x"5472802e",
  1184 => x"80c43873",
  1185 => x"80dcc00b",
  1186 => x"80d7d80c",
  1187 => x"80d5ec53",
  1188 => x"80dcbc52",
  1189 => x"5ea3952d",
  1190 => x"ff177052",
  1191 => x"53a2e42d",
  1192 => x"72882c51",
  1193 => x"a2e42da0",
  1194 => x"51a2af2d",
  1195 => x"7951a2e4",
  1196 => x"2da051a2",
  1197 => x"af2d7a51",
  1198 => x"a2e42d80",
  1199 => x"dcbc5280",
  1200 => x"dbf851a3",
  1201 => x"952dff19",
  1202 => x"59788025",
  1203 => x"ff8338a5",
  1204 => x"da0480db",
  1205 => x"d0085884",
  1206 => x"805680db",
  1207 => x"ec5180cd",
  1208 => x"8a2dfc80",
  1209 => x"16811656",
  1210 => x"56a48a04",
  1211 => x"80dbf008",
  1212 => x"f80c7d8a",
  1213 => x"387f5280",
  1214 => x"dbf851a3",
  1215 => x"952d8051",
  1216 => x"86da2d77",
  1217 => x"802e8838",
  1218 => x"80d7dc51",
  1219 => x"a6930480",
  1220 => x"d99c51af",
  1221 => x"982d7780",
  1222 => x"dbd00c02",
  1223 => x"80c0050d",
  1224 => x"0402ec05",
  1225 => x"0d80dcbc",
  1226 => x"0b80d7d8",
  1227 => x"0c80dcbc",
  1228 => x"55807581",
  1229 => x"b72d80d9",
  1230 => x"c00851a2",
  1231 => x"e42dba51",
  1232 => x"a2af2dff",
  1233 => x"b8087098",
  1234 => x"2a5254a2",
  1235 => x"e42d7390",
  1236 => x"2a7081ff",
  1237 => x"065253a2",
  1238 => x"e42d7388",
  1239 => x"2a7081ff",
  1240 => x"065253a2",
  1241 => x"e42d7381",
  1242 => x"ff0651a2",
  1243 => x"e42d7452",
  1244 => x"80dbf851",
  1245 => x"a3952d80",
  1246 => x"d7dc51af",
  1247 => x"982d80d9",
  1248 => x"c0088405",
  1249 => x"80d9c00c",
  1250 => x"0294050d",
  1251 => x"04800b80",
  1252 => x"d9c00c04",
  1253 => x"02ec050d",
  1254 => x"840bec0c",
  1255 => x"acd52da9",
  1256 => x"8a2d81f9",
  1257 => x"2d8353ac",
  1258 => x"b82d8151",
  1259 => x"858d2dff",
  1260 => x"13537280",
  1261 => x"25f13884",
  1262 => x"0bec0c80",
  1263 => x"d5f45186",
  1264 => x"a02d80c1",
  1265 => x"922d80db",
  1266 => x"d008802e",
  1267 => x"81a538a3",
  1268 => x"bc5180d4",
  1269 => x"902d80d6",
  1270 => x"8c5280db",
  1271 => x"f851a395",
  1272 => x"2d80d7dc",
  1273 => x"51af982d",
  1274 => x"acf72da9",
  1275 => x"962dafab",
  1276 => x"2d80d7f0",
  1277 => x"0b80f52d",
  1278 => x"80da8c08",
  1279 => x"70810655",
  1280 => x"56547280",
  1281 => x"2e853873",
  1282 => x"84075474",
  1283 => x"812a7081",
  1284 => x"06515372",
  1285 => x"802e8538",
  1286 => x"73820754",
  1287 => x"74822a70",
  1288 => x"81065153",
  1289 => x"72802e85",
  1290 => x"38738107",
  1291 => x"5474832a",
  1292 => x"70810651",
  1293 => x"5372802e",
  1294 => x"85387388",
  1295 => x"07547484",
  1296 => x"2a708106",
  1297 => x"51537280",
  1298 => x"2e853873",
  1299 => x"90075474",
  1300 => x"852a7081",
  1301 => x"06515372",
  1302 => x"802e8538",
  1303 => x"73a00754",
  1304 => x"73fc0c86",
  1305 => x"5380dbd0",
  1306 => x"08833884",
  1307 => x"5372ec0c",
  1308 => x"a7eb0480",
  1309 => x"0b80dbd0",
  1310 => x"0c029405",
  1311 => x"0d047198",
  1312 => x"0c04ffb0",
  1313 => x"0880dbd0",
  1314 => x"0c04810b",
  1315 => x"ffb00c04",
  1316 => x"800bffb0",
  1317 => x"0c0402f4",
  1318 => x"050daaa4",
  1319 => x"0480dbd0",
  1320 => x"0881f02e",
  1321 => x"0981068a",
  1322 => x"38810b80",
  1323 => x"da840caa",
  1324 => x"a40480db",
  1325 => x"d00881e0",
  1326 => x"2e098106",
  1327 => x"8a38810b",
  1328 => x"80da880c",
  1329 => x"aaa40480",
  1330 => x"dbd00852",
  1331 => x"80da8808",
  1332 => x"802e8938",
  1333 => x"80dbd008",
  1334 => x"81800552",
  1335 => x"71842c72",
  1336 => x"8f065353",
  1337 => x"80da8408",
  1338 => x"802e9a38",
  1339 => x"72842980",
  1340 => x"d9c40572",
  1341 => x"1381712b",
  1342 => x"70097308",
  1343 => x"06730c51",
  1344 => x"5353aa98",
  1345 => x"04728429",
  1346 => x"80d9c405",
  1347 => x"72138371",
  1348 => x"2b720807",
  1349 => x"720c5353",
  1350 => x"800b80da",
  1351 => x"880c800b",
  1352 => x"80da840c",
  1353 => x"80dd8051",
  1354 => x"abab2d80",
  1355 => x"dbd008ff",
  1356 => x"24feea38",
  1357 => x"800b80db",
  1358 => x"d00c028c",
  1359 => x"050d0402",
  1360 => x"f8050d80",
  1361 => x"d9c4528f",
  1362 => x"51807270",
  1363 => x"8405540c",
  1364 => x"ff115170",
  1365 => x"8025f238",
  1366 => x"0288050d",
  1367 => x"0402f005",
  1368 => x"0d7551a9",
  1369 => x"902d7082",
  1370 => x"2cfc0680",
  1371 => x"d9c41172",
  1372 => x"109e0671",
  1373 => x"0870722a",
  1374 => x"70830682",
  1375 => x"742b7009",
  1376 => x"7406760c",
  1377 => x"54515657",
  1378 => x"535153a9",
  1379 => x"8a2d7180",
  1380 => x"dbd00c02",
  1381 => x"90050d04",
  1382 => x"02fc050d",
  1383 => x"72518071",
  1384 => x"0c800b84",
  1385 => x"120c0284",
  1386 => x"050d0402",
  1387 => x"f0050d75",
  1388 => x"70088412",
  1389 => x"08535353",
  1390 => x"ff547171",
  1391 => x"2ea838a9",
  1392 => x"902d8413",
  1393 => x"08708429",
  1394 => x"14881170",
  1395 => x"087081ff",
  1396 => x"06841808",
  1397 => x"81118706",
  1398 => x"841a0c53",
  1399 => x"51555151",
  1400 => x"51a98a2d",
  1401 => x"71547380",
  1402 => x"dbd00c02",
  1403 => x"90050d04",
  1404 => x"02f8050d",
  1405 => x"a9902de0",
  1406 => x"08708b2a",
  1407 => x"70810651",
  1408 => x"52527080",
  1409 => x"2ea13880",
  1410 => x"dd800870",
  1411 => x"842980dd",
  1412 => x"88057381",
  1413 => x"ff06710c",
  1414 => x"515180dd",
  1415 => x"80088111",
  1416 => x"870680dd",
  1417 => x"800c5180",
  1418 => x"0b80dda8",
  1419 => x"0ca9822d",
  1420 => x"a98a2d02",
  1421 => x"88050d04",
  1422 => x"02fc050d",
  1423 => x"a9902d81",
  1424 => x"0b80dda8",
  1425 => x"0ca98a2d",
  1426 => x"80dda808",
  1427 => x"5170f938",
  1428 => x"0284050d",
  1429 => x"0402fc05",
  1430 => x"0d80dd80",
  1431 => x"51ab982d",
  1432 => x"aabf2dab",
  1433 => x"f051a8fe",
  1434 => x"2d028405",
  1435 => x"0d0480dd",
  1436 => x"b40880db",
  1437 => x"d00c0402",
  1438 => x"fc050d81",
  1439 => x"0b80da90",
  1440 => x"0c815185",
  1441 => x"8d2d0284",
  1442 => x"050d0402",
  1443 => x"fc050dad",
  1444 => x"9504a996",
  1445 => x"2d80f651",
  1446 => x"aadd2d80",
  1447 => x"dbd008f2",
  1448 => x"3880da51",
  1449 => x"aadd2d80",
  1450 => x"dbd008e6",
  1451 => x"3880dbd0",
  1452 => x"0880da90",
  1453 => x"0c80dbd0",
  1454 => x"0851858d",
  1455 => x"2d028405",
  1456 => x"0d0402ec",
  1457 => x"050d7654",
  1458 => x"8052870b",
  1459 => x"881580f5",
  1460 => x"2d565374",
  1461 => x"72248338",
  1462 => x"a0537251",
  1463 => x"83842d81",
  1464 => x"128b1580",
  1465 => x"f52d5452",
  1466 => x"727225de",
  1467 => x"38029405",
  1468 => x"0d0402f0",
  1469 => x"050d80dd",
  1470 => x"b4085481",
  1471 => x"f92d800b",
  1472 => x"80ddb80c",
  1473 => x"7308802e",
  1474 => x"81893882",
  1475 => x"0b80dbe4",
  1476 => x"0c80ddb8",
  1477 => x"088f0680",
  1478 => x"dbe00c73",
  1479 => x"08527183",
  1480 => x"2e963871",
  1481 => x"83268938",
  1482 => x"71812eb0",
  1483 => x"38aefc04",
  1484 => x"71852ea0",
  1485 => x"38aefc04",
  1486 => x"881480f5",
  1487 => x"2d841508",
  1488 => x"80d69c53",
  1489 => x"545286a0",
  1490 => x"2d718429",
  1491 => x"13700852",
  1492 => x"52af8004",
  1493 => x"7351adc2",
  1494 => x"2daefc04",
  1495 => x"80da8c08",
  1496 => x"8815082c",
  1497 => x"70810651",
  1498 => x"5271802e",
  1499 => x"883880d6",
  1500 => x"a051aef9",
  1501 => x"0480d6a4",
  1502 => x"5186a02d",
  1503 => x"84140851",
  1504 => x"86a02d80",
  1505 => x"ddb80881",
  1506 => x"0580ddb8",
  1507 => x"0c8c1454",
  1508 => x"ae840402",
  1509 => x"90050d04",
  1510 => x"7180ddb4",
  1511 => x"0cadf22d",
  1512 => x"80ddb808",
  1513 => x"ff0580dd",
  1514 => x"bc0c0402",
  1515 => x"e8050d80",
  1516 => x"ddb40880",
  1517 => x"ddc00857",
  1518 => x"5580f651",
  1519 => x"aadd2d80",
  1520 => x"dbd00881",
  1521 => x"2a708106",
  1522 => x"51527180",
  1523 => x"2ea438af",
  1524 => x"d504a996",
  1525 => x"2d80f651",
  1526 => x"aadd2d80",
  1527 => x"dbd008f2",
  1528 => x"3880da90",
  1529 => x"08813270",
  1530 => x"80da900c",
  1531 => x"70525285",
  1532 => x"8d2d800b",
  1533 => x"80ddac0c",
  1534 => x"800b80dd",
  1535 => x"b00c80da",
  1536 => x"9008838d",
  1537 => x"3880da51",
  1538 => x"aadd2d80",
  1539 => x"dbd00880",
  1540 => x"2e8c3880",
  1541 => x"ddac0881",
  1542 => x"800780dd",
  1543 => x"ac0c80d9",
  1544 => x"51aadd2d",
  1545 => x"80dbd008",
  1546 => x"802e8c38",
  1547 => x"80ddac08",
  1548 => x"80c00780",
  1549 => x"ddac0c81",
  1550 => x"9451aadd",
  1551 => x"2d80dbd0",
  1552 => x"08802e8b",
  1553 => x"3880ddac",
  1554 => x"08900780",
  1555 => x"ddac0c81",
  1556 => x"9151aadd",
  1557 => x"2d80dbd0",
  1558 => x"08802e8b",
  1559 => x"3880ddac",
  1560 => x"08a00780",
  1561 => x"ddac0c81",
  1562 => x"f551aadd",
  1563 => x"2d80dbd0",
  1564 => x"08802e8b",
  1565 => x"3880ddac",
  1566 => x"08810780",
  1567 => x"ddac0c81",
  1568 => x"f251aadd",
  1569 => x"2d80dbd0",
  1570 => x"08802e8b",
  1571 => x"3880ddac",
  1572 => x"08820780",
  1573 => x"ddac0c81",
  1574 => x"eb51aadd",
  1575 => x"2d80dbd0",
  1576 => x"08802e8b",
  1577 => x"3880ddac",
  1578 => x"08840780",
  1579 => x"ddac0c81",
  1580 => x"f451aadd",
  1581 => x"2d80dbd0",
  1582 => x"08802e8b",
  1583 => x"3880ddac",
  1584 => x"08880780",
  1585 => x"ddac0c80",
  1586 => x"d851aadd",
  1587 => x"2d80dbd0",
  1588 => x"08802e8c",
  1589 => x"3880ddb0",
  1590 => x"08818007",
  1591 => x"80ddb00c",
  1592 => x"9251aadd",
  1593 => x"2d80dbd0",
  1594 => x"08802e8c",
  1595 => x"3880ddb0",
  1596 => x"0880c007",
  1597 => x"80ddb00c",
  1598 => x"9451aadd",
  1599 => x"2d80dbd0",
  1600 => x"08802e8b",
  1601 => x"3880ddb0",
  1602 => x"08900780",
  1603 => x"ddb00c91",
  1604 => x"51aadd2d",
  1605 => x"80dbd008",
  1606 => x"802e8b38",
  1607 => x"80ddb008",
  1608 => x"a00780dd",
  1609 => x"b00c9d51",
  1610 => x"aadd2d80",
  1611 => x"dbd00880",
  1612 => x"2e8b3880",
  1613 => x"ddb00881",
  1614 => x"0780ddb0",
  1615 => x"0c9b51aa",
  1616 => x"dd2d80db",
  1617 => x"d008802e",
  1618 => x"8b3880dd",
  1619 => x"b0088207",
  1620 => x"80ddb00c",
  1621 => x"9c51aadd",
  1622 => x"2d80dbd0",
  1623 => x"08802e8b",
  1624 => x"3880ddb0",
  1625 => x"08840780",
  1626 => x"ddb00ca3",
  1627 => x"51aadd2d",
  1628 => x"80dbd008",
  1629 => x"802e8b38",
  1630 => x"80ddb008",
  1631 => x"880780dd",
  1632 => x"b00c81fd",
  1633 => x"51aadd2d",
  1634 => x"81fa51aa",
  1635 => x"dd2db8e6",
  1636 => x"0481f551",
  1637 => x"aadd2d80",
  1638 => x"dbd00881",
  1639 => x"2a708106",
  1640 => x"51527180",
  1641 => x"2eb33880",
  1642 => x"ddbc0852",
  1643 => x"71802e8a",
  1644 => x"38ff1280",
  1645 => x"ddbc0cb3",
  1646 => x"d90480dd",
  1647 => x"b8081080",
  1648 => x"ddb80805",
  1649 => x"70842916",
  1650 => x"51528812",
  1651 => x"08802e89",
  1652 => x"38ff5188",
  1653 => x"12085271",
  1654 => x"2d81f251",
  1655 => x"aadd2d80",
  1656 => x"dbd00881",
  1657 => x"2a708106",
  1658 => x"51527180",
  1659 => x"2eb43880",
  1660 => x"ddb808ff",
  1661 => x"1180ddbc",
  1662 => x"08565353",
  1663 => x"7372258a",
  1664 => x"38811480",
  1665 => x"ddbc0cb4",
  1666 => x"a2047210",
  1667 => x"13708429",
  1668 => x"16515288",
  1669 => x"1208802e",
  1670 => x"8938fe51",
  1671 => x"88120852",
  1672 => x"712d81fd",
  1673 => x"51aadd2d",
  1674 => x"80dbd008",
  1675 => x"812a7081",
  1676 => x"06515271",
  1677 => x"802eb138",
  1678 => x"80ddbc08",
  1679 => x"802e8a38",
  1680 => x"800b80dd",
  1681 => x"bc0cb4e8",
  1682 => x"0480ddb8",
  1683 => x"081080dd",
  1684 => x"b8080570",
  1685 => x"84291651",
  1686 => x"52881208",
  1687 => x"802e8938",
  1688 => x"fd518812",
  1689 => x"0852712d",
  1690 => x"81fa51aa",
  1691 => x"dd2d80db",
  1692 => x"d008812a",
  1693 => x"70810651",
  1694 => x"5271802e",
  1695 => x"b13880dd",
  1696 => x"b808ff11",
  1697 => x"545280dd",
  1698 => x"bc087325",
  1699 => x"89387280",
  1700 => x"ddbc0cb5",
  1701 => x"ae047110",
  1702 => x"12708429",
  1703 => x"16515288",
  1704 => x"1208802e",
  1705 => x"8938fc51",
  1706 => x"88120852",
  1707 => x"712d80dd",
  1708 => x"bc087053",
  1709 => x"5473802e",
  1710 => x"8a388c15",
  1711 => x"ff155555",
  1712 => x"b5b50482",
  1713 => x"0b80dbe4",
  1714 => x"0c718f06",
  1715 => x"80dbe00c",
  1716 => x"81eb51aa",
  1717 => x"dd2d80db",
  1718 => x"d008812a",
  1719 => x"70810651",
  1720 => x"5271802e",
  1721 => x"ad387408",
  1722 => x"852e0981",
  1723 => x"06a43888",
  1724 => x"1580f52d",
  1725 => x"ff055271",
  1726 => x"881681b7",
  1727 => x"2d71982b",
  1728 => x"52718025",
  1729 => x"8838800b",
  1730 => x"881681b7",
  1731 => x"2d7451ad",
  1732 => x"c22d81f4",
  1733 => x"51aadd2d",
  1734 => x"80dbd008",
  1735 => x"812a7081",
  1736 => x"06515271",
  1737 => x"802eb338",
  1738 => x"7408852e",
  1739 => x"098106aa",
  1740 => x"38881580",
  1741 => x"f52d8105",
  1742 => x"52718816",
  1743 => x"81b72d71",
  1744 => x"81ff068b",
  1745 => x"1680f52d",
  1746 => x"54527272",
  1747 => x"27873872",
  1748 => x"881681b7",
  1749 => x"2d7451ad",
  1750 => x"c22d80da",
  1751 => x"51aadd2d",
  1752 => x"80dbd008",
  1753 => x"812a7081",
  1754 => x"06515271",
  1755 => x"802e81ad",
  1756 => x"3880ddb4",
  1757 => x"0880ddbc",
  1758 => x"08555373",
  1759 => x"802e8a38",
  1760 => x"8c13ff15",
  1761 => x"5553b6fb",
  1762 => x"04720852",
  1763 => x"71822ea6",
  1764 => x"38718226",
  1765 => x"89387181",
  1766 => x"2eaa38b8",
  1767 => x"9d047183",
  1768 => x"2eb43871",
  1769 => x"842e0981",
  1770 => x"0680f238",
  1771 => x"88130851",
  1772 => x"af982db8",
  1773 => x"9d0480dd",
  1774 => x"bc085188",
  1775 => x"13085271",
  1776 => x"2db89d04",
  1777 => x"810b8814",
  1778 => x"082b80da",
  1779 => x"8c083280",
  1780 => x"da8c0cb7",
  1781 => x"f1048813",
  1782 => x"80f52d81",
  1783 => x"058b1480",
  1784 => x"f52d5354",
  1785 => x"71742483",
  1786 => x"38805473",
  1787 => x"881481b7",
  1788 => x"2dadf22d",
  1789 => x"b89d0475",
  1790 => x"08802ea4",
  1791 => x"38750851",
  1792 => x"aadd2d80",
  1793 => x"dbd00881",
  1794 => x"06527180",
  1795 => x"2e8c3880",
  1796 => x"ddbc0851",
  1797 => x"84160852",
  1798 => x"712d8816",
  1799 => x"5675d838",
  1800 => x"8054800b",
  1801 => x"80dbe40c",
  1802 => x"738f0680",
  1803 => x"dbe00ca0",
  1804 => x"527380dd",
  1805 => x"bc082e09",
  1806 => x"81069938",
  1807 => x"80ddb808",
  1808 => x"ff057432",
  1809 => x"70098105",
  1810 => x"7072079f",
  1811 => x"2a917131",
  1812 => x"51515353",
  1813 => x"71518384",
  1814 => x"2d811454",
  1815 => x"8e7425c2",
  1816 => x"3880da90",
  1817 => x"08527180",
  1818 => x"dbd00c02",
  1819 => x"98050d04",
  1820 => x"02f4050d",
  1821 => x"d45281ff",
  1822 => x"720c7108",
  1823 => x"5381ff72",
  1824 => x"0c72882b",
  1825 => x"83fe8006",
  1826 => x"72087081",
  1827 => x"ff065152",
  1828 => x"5381ff72",
  1829 => x"0c727107",
  1830 => x"882b7208",
  1831 => x"7081ff06",
  1832 => x"51525381",
  1833 => x"ff720c72",
  1834 => x"7107882b",
  1835 => x"72087081",
  1836 => x"ff067207",
  1837 => x"80dbd00c",
  1838 => x"5253028c",
  1839 => x"050d0402",
  1840 => x"f4050d74",
  1841 => x"767181ff",
  1842 => x"06d40c53",
  1843 => x"5380ddc4",
  1844 => x"08853871",
  1845 => x"892b5271",
  1846 => x"982ad40c",
  1847 => x"71902a70",
  1848 => x"81ff06d4",
  1849 => x"0c517188",
  1850 => x"2a7081ff",
  1851 => x"06d40c51",
  1852 => x"7181ff06",
  1853 => x"d40c7290",
  1854 => x"2a7081ff",
  1855 => x"06d40c51",
  1856 => x"d4087081",
  1857 => x"ff065151",
  1858 => x"82b8bf52",
  1859 => x"7081ff2e",
  1860 => x"09810694",
  1861 => x"3881ff0b",
  1862 => x"d40cd408",
  1863 => x"7081ff06",
  1864 => x"ff145451",
  1865 => x"5171e538",
  1866 => x"7080dbd0",
  1867 => x"0c028c05",
  1868 => x"0d0402fc",
  1869 => x"050d81c7",
  1870 => x"5181ff0b",
  1871 => x"d40cff11",
  1872 => x"51708025",
  1873 => x"f4380284",
  1874 => x"050d0402",
  1875 => x"f4050d81",
  1876 => x"ff0bd40c",
  1877 => x"93538052",
  1878 => x"87fc80c1",
  1879 => x"51b9bf2d",
  1880 => x"80dbd008",
  1881 => x"8b3881ff",
  1882 => x"0bd40c81",
  1883 => x"53baf904",
  1884 => x"bab22dff",
  1885 => x"135372de",
  1886 => x"387280db",
  1887 => x"d00c028c",
  1888 => x"050d0402",
  1889 => x"ec050d81",
  1890 => x"0b80ddc4",
  1891 => x"0c8454d0",
  1892 => x"08708f2a",
  1893 => x"70810651",
  1894 => x"515372f3",
  1895 => x"3872d00c",
  1896 => x"bab22d80",
  1897 => x"d6a85186",
  1898 => x"a02dd008",
  1899 => x"708f2a70",
  1900 => x"81065151",
  1901 => x"5372f338",
  1902 => x"810bd00c",
  1903 => x"b1538052",
  1904 => x"84d480c0",
  1905 => x"51b9bf2d",
  1906 => x"80dbd008",
  1907 => x"812e9338",
  1908 => x"72822ebf",
  1909 => x"38ff1353",
  1910 => x"72e438ff",
  1911 => x"145473ff",
  1912 => x"ae38bab2",
  1913 => x"2d83aa52",
  1914 => x"849c80c8",
  1915 => x"51b9bf2d",
  1916 => x"80dbd008",
  1917 => x"812e0981",
  1918 => x"069338b8",
  1919 => x"f02d80db",
  1920 => x"d00883ff",
  1921 => x"ff065372",
  1922 => x"83aa2e9f",
  1923 => x"38bacb2d",
  1924 => x"bca60480",
  1925 => x"d6b45186",
  1926 => x"a02d8053",
  1927 => x"bdfb0480",
  1928 => x"d6cc5186",
  1929 => x"a02d8054",
  1930 => x"bdcc0481",
  1931 => x"ff0bd40c",
  1932 => x"b154bab2",
  1933 => x"2d8fcf53",
  1934 => x"805287fc",
  1935 => x"80f751b9",
  1936 => x"bf2d80db",
  1937 => x"d0085580",
  1938 => x"dbd00881",
  1939 => x"2e098106",
  1940 => x"9c3881ff",
  1941 => x"0bd40c82",
  1942 => x"0a52849c",
  1943 => x"80e951b9",
  1944 => x"bf2d80db",
  1945 => x"d008802e",
  1946 => x"8d38bab2",
  1947 => x"2dff1353",
  1948 => x"72c638bd",
  1949 => x"bf0481ff",
  1950 => x"0bd40c80",
  1951 => x"dbd00852",
  1952 => x"87fc80fa",
  1953 => x"51b9bf2d",
  1954 => x"80dbd008",
  1955 => x"b23881ff",
  1956 => x"0bd40cd4",
  1957 => x"085381ff",
  1958 => x"0bd40c81",
  1959 => x"ff0bd40c",
  1960 => x"81ff0bd4",
  1961 => x"0c81ff0b",
  1962 => x"d40c7286",
  1963 => x"2a708106",
  1964 => x"76565153",
  1965 => x"72963880",
  1966 => x"dbd00854",
  1967 => x"bdcc0473",
  1968 => x"822efedb",
  1969 => x"38ff1454",
  1970 => x"73fee738",
  1971 => x"7380ddc4",
  1972 => x"0c738b38",
  1973 => x"815287fc",
  1974 => x"80d051b9",
  1975 => x"bf2d81ff",
  1976 => x"0bd40cd0",
  1977 => x"08708f2a",
  1978 => x"70810651",
  1979 => x"515372f3",
  1980 => x"3872d00c",
  1981 => x"81ff0bd4",
  1982 => x"0c815372",
  1983 => x"80dbd00c",
  1984 => x"0294050d",
  1985 => x"0402e805",
  1986 => x"0d785580",
  1987 => x"5681ff0b",
  1988 => x"d40cd008",
  1989 => x"708f2a70",
  1990 => x"81065151",
  1991 => x"5372f338",
  1992 => x"82810bd0",
  1993 => x"0c81ff0b",
  1994 => x"d40c7752",
  1995 => x"87fc80d1",
  1996 => x"51b9bf2d",
  1997 => x"80dbc6df",
  1998 => x"5480dbd0",
  1999 => x"08802e8b",
  2000 => x"3880d6ec",
  2001 => x"5186a02d",
  2002 => x"bf9f0481",
  2003 => x"ff0bd40c",
  2004 => x"d4087081",
  2005 => x"ff065153",
  2006 => x"7281fe2e",
  2007 => x"0981069e",
  2008 => x"3880ff53",
  2009 => x"b8f02d80",
  2010 => x"dbd00875",
  2011 => x"70840557",
  2012 => x"0cff1353",
  2013 => x"728025ec",
  2014 => x"388156bf",
  2015 => x"8404ff14",
  2016 => x"5473c838",
  2017 => x"81ff0bd4",
  2018 => x"0c81ff0b",
  2019 => x"d40cd008",
  2020 => x"708f2a70",
  2021 => x"81065151",
  2022 => x"5372f338",
  2023 => x"72d00c75",
  2024 => x"80dbd00c",
  2025 => x"0298050d",
  2026 => x"0402e805",
  2027 => x"0d77797b",
  2028 => x"58555580",
  2029 => x"53727625",
  2030 => x"a3387470",
  2031 => x"81055680",
  2032 => x"f52d7470",
  2033 => x"81055680",
  2034 => x"f52d5252",
  2035 => x"71712e86",
  2036 => x"388151bf",
  2037 => x"de048113",
  2038 => x"53bfb504",
  2039 => x"80517080",
  2040 => x"dbd00c02",
  2041 => x"98050d04",
  2042 => x"02ec050d",
  2043 => x"76557480",
  2044 => x"2e80c438",
  2045 => x"9a1580e0",
  2046 => x"2d5180ce",
  2047 => x"952d80db",
  2048 => x"d00880db",
  2049 => x"d00880e3",
  2050 => x"f80c80db",
  2051 => x"d0085454",
  2052 => x"80e3d408",
  2053 => x"802e9b38",
  2054 => x"941580e0",
  2055 => x"2d5180ce",
  2056 => x"952d80db",
  2057 => x"d008902b",
  2058 => x"83fff00a",
  2059 => x"06707507",
  2060 => x"51537280",
  2061 => x"e3f80c80",
  2062 => x"e3f80853",
  2063 => x"72802e9e",
  2064 => x"3880e3cc",
  2065 => x"08fe1471",
  2066 => x"2980e3e0",
  2067 => x"080580e3",
  2068 => x"fc0c7084",
  2069 => x"2b80e3d8",
  2070 => x"0c5480c1",
  2071 => x"8d0480e3",
  2072 => x"e40880e3",
  2073 => x"f80c80e3",
  2074 => x"e80880e3",
  2075 => x"fc0c80e3",
  2076 => x"d408802e",
  2077 => x"8c3880e3",
  2078 => x"cc08842b",
  2079 => x"5380c188",
  2080 => x"0480e3ec",
  2081 => x"08842b53",
  2082 => x"7280e3d8",
  2083 => x"0c029405",
  2084 => x"0d0402d8",
  2085 => x"050d800b",
  2086 => x"80e3d40c",
  2087 => x"8454bb83",
  2088 => x"2d80dbd0",
  2089 => x"08802e98",
  2090 => x"3880ddc8",
  2091 => x"528051be",
  2092 => x"852d80db",
  2093 => x"d008802e",
  2094 => x"8738fe54",
  2095 => x"80c1c804",
  2096 => x"ff145473",
  2097 => x"8024d738",
  2098 => x"738e3880",
  2099 => x"d6fc5186",
  2100 => x"a02d7355",
  2101 => x"80c7a504",
  2102 => x"8056810b",
  2103 => x"80e4800c",
  2104 => x"885380d7",
  2105 => x"905280dd",
  2106 => x"fe51bfa9",
  2107 => x"2d80dbd0",
  2108 => x"08762e09",
  2109 => x"81068938",
  2110 => x"80dbd008",
  2111 => x"80e4800c",
  2112 => x"885380d7",
  2113 => x"9c5280de",
  2114 => x"9a51bfa9",
  2115 => x"2d80dbd0",
  2116 => x"08893880",
  2117 => x"dbd00880",
  2118 => x"e4800c80",
  2119 => x"e4800880",
  2120 => x"2e818438",
  2121 => x"80e18e0b",
  2122 => x"80f52d80",
  2123 => x"e18f0b80",
  2124 => x"f52d7198",
  2125 => x"2b71902b",
  2126 => x"0780e190",
  2127 => x"0b80f52d",
  2128 => x"70882b72",
  2129 => x"0780e191",
  2130 => x"0b80f52d",
  2131 => x"710780e1",
  2132 => x"c60b80f5",
  2133 => x"2d80e1c7",
  2134 => x"0b80f52d",
  2135 => x"71882b07",
  2136 => x"535f5452",
  2137 => x"5a565755",
  2138 => x"7381abaa",
  2139 => x"2e098106",
  2140 => x"90387551",
  2141 => x"80cde42d",
  2142 => x"80dbd008",
  2143 => x"5680c390",
  2144 => x"047382d4",
  2145 => x"d52e8938",
  2146 => x"80d7a851",
  2147 => x"80c3dd04",
  2148 => x"80ddc852",
  2149 => x"7551be85",
  2150 => x"2d80dbd0",
  2151 => x"085580db",
  2152 => x"d008802e",
  2153 => x"83ff3888",
  2154 => x"5380d79c",
  2155 => x"5280de9a",
  2156 => x"51bfa92d",
  2157 => x"80dbd008",
  2158 => x"8b38810b",
  2159 => x"80e3d40c",
  2160 => x"80c3e404",
  2161 => x"885380d7",
  2162 => x"905280dd",
  2163 => x"fe51bfa9",
  2164 => x"2d80dbd0",
  2165 => x"08802e8c",
  2166 => x"3880d7bc",
  2167 => x"5186a02d",
  2168 => x"80c4c304",
  2169 => x"80e1c60b",
  2170 => x"80f52d54",
  2171 => x"7380d52e",
  2172 => x"09810680",
  2173 => x"ce3880e1",
  2174 => x"c70b80f5",
  2175 => x"2d547381",
  2176 => x"aa2e0981",
  2177 => x"06bd3880",
  2178 => x"0b80ddc8",
  2179 => x"0b80f52d",
  2180 => x"56547481",
  2181 => x"e92e8338",
  2182 => x"81547481",
  2183 => x"eb2e8c38",
  2184 => x"80557375",
  2185 => x"2e098106",
  2186 => x"82fb3880",
  2187 => x"ddd30b80",
  2188 => x"f52d5574",
  2189 => x"8e3880dd",
  2190 => x"d40b80f5",
  2191 => x"2d547382",
  2192 => x"2e873880",
  2193 => x"5580c7a5",
  2194 => x"0480ddd5",
  2195 => x"0b80f52d",
  2196 => x"7080e3cc",
  2197 => x"0cff0580",
  2198 => x"e3d00c80",
  2199 => x"ddd60b80",
  2200 => x"f52d80dd",
  2201 => x"d70b80f5",
  2202 => x"2d587605",
  2203 => x"77828029",
  2204 => x"057080e3",
  2205 => x"dc0c80dd",
  2206 => x"d80b80f5",
  2207 => x"2d7080e3",
  2208 => x"f00c80e3",
  2209 => x"d4085957",
  2210 => x"5876802e",
  2211 => x"81b83888",
  2212 => x"5380d79c",
  2213 => x"5280de9a",
  2214 => x"51bfa92d",
  2215 => x"80dbd008",
  2216 => x"82833880",
  2217 => x"e3cc0870",
  2218 => x"842b80e3",
  2219 => x"d80c7080",
  2220 => x"e3ec0c80",
  2221 => x"dded0b80",
  2222 => x"f52d80dd",
  2223 => x"ec0b80f5",
  2224 => x"2d718280",
  2225 => x"290580dd",
  2226 => x"ee0b80f5",
  2227 => x"2d708480",
  2228 => x"80291280",
  2229 => x"ddef0b80",
  2230 => x"f52d7081",
  2231 => x"800a2912",
  2232 => x"7080e3f4",
  2233 => x"0c80e3f0",
  2234 => x"08712980",
  2235 => x"e3dc0805",
  2236 => x"7080e3e0",
  2237 => x"0c80ddf5",
  2238 => x"0b80f52d",
  2239 => x"80ddf40b",
  2240 => x"80f52d71",
  2241 => x"82802905",
  2242 => x"80ddf60b",
  2243 => x"80f52d70",
  2244 => x"84808029",
  2245 => x"1280ddf7",
  2246 => x"0b80f52d",
  2247 => x"70982b81",
  2248 => x"f00a0672",
  2249 => x"057080e3",
  2250 => x"e40cfe11",
  2251 => x"7e297705",
  2252 => x"80e3e80c",
  2253 => x"52595243",
  2254 => x"545e5152",
  2255 => x"59525d57",
  2256 => x"595780c7",
  2257 => x"9e0480dd",
  2258 => x"da0b80f5",
  2259 => x"2d80ddd9",
  2260 => x"0b80f52d",
  2261 => x"71828029",
  2262 => x"057080e3",
  2263 => x"d80c70a0",
  2264 => x"2983ff05",
  2265 => x"70892a70",
  2266 => x"80e3ec0c",
  2267 => x"80dddf0b",
  2268 => x"80f52d80",
  2269 => x"ddde0b80",
  2270 => x"f52d7182",
  2271 => x"80290570",
  2272 => x"80e3f40c",
  2273 => x"7b71291e",
  2274 => x"7080e3e8",
  2275 => x"0c7d80e3",
  2276 => x"e40c7305",
  2277 => x"80e3e00c",
  2278 => x"555e5151",
  2279 => x"55558051",
  2280 => x"bfe82d81",
  2281 => x"557480db",
  2282 => x"d00c02a8",
  2283 => x"050d0402",
  2284 => x"ec050d76",
  2285 => x"70872c71",
  2286 => x"80ff0655",
  2287 => x"565480e3",
  2288 => x"d4088a38",
  2289 => x"73882c74",
  2290 => x"81ff0654",
  2291 => x"5580ddc8",
  2292 => x"5280e3dc",
  2293 => x"081551be",
  2294 => x"852d80db",
  2295 => x"d0085480",
  2296 => x"dbd00880",
  2297 => x"2ebb3880",
  2298 => x"e3d40880",
  2299 => x"2e9c3872",
  2300 => x"842980dd",
  2301 => x"c8057008",
  2302 => x"525380cd",
  2303 => x"e42d80db",
  2304 => x"d008f00a",
  2305 => x"065380c8",
  2306 => x"9f047210",
  2307 => x"80ddc805",
  2308 => x"7080e02d",
  2309 => x"525380ce",
  2310 => x"952d80db",
  2311 => x"d0085372",
  2312 => x"547380db",
  2313 => x"d00c0294",
  2314 => x"050d0402",
  2315 => x"e0050d79",
  2316 => x"70842c80",
  2317 => x"e3fc0805",
  2318 => x"718f0652",
  2319 => x"5553728a",
  2320 => x"3880ddc8",
  2321 => x"527351be",
  2322 => x"852d72a0",
  2323 => x"2980ddc8",
  2324 => x"05548074",
  2325 => x"80f52d56",
  2326 => x"5374732e",
  2327 => x"83388153",
  2328 => x"7481e52e",
  2329 => x"81f53881",
  2330 => x"70740654",
  2331 => x"5872802e",
  2332 => x"81e9388b",
  2333 => x"1480f52d",
  2334 => x"70832a79",
  2335 => x"06585676",
  2336 => x"9c3880da",
  2337 => x"94085372",
  2338 => x"89387280",
  2339 => x"e1c80b81",
  2340 => x"b72d7680",
  2341 => x"da940c73",
  2342 => x"5380cadd",
  2343 => x"04758f2e",
  2344 => x"09810681",
  2345 => x"b638749f",
  2346 => x"068d2980",
  2347 => x"e1bb1151",
  2348 => x"53811480",
  2349 => x"f52d7370",
  2350 => x"81055581",
  2351 => x"b72d8314",
  2352 => x"80f52d73",
  2353 => x"70810555",
  2354 => x"81b72d85",
  2355 => x"1480f52d",
  2356 => x"73708105",
  2357 => x"5581b72d",
  2358 => x"871480f5",
  2359 => x"2d737081",
  2360 => x"055581b7",
  2361 => x"2d891480",
  2362 => x"f52d7370",
  2363 => x"81055581",
  2364 => x"b72d8e14",
  2365 => x"80f52d73",
  2366 => x"70810555",
  2367 => x"81b72d90",
  2368 => x"1480f52d",
  2369 => x"73708105",
  2370 => x"5581b72d",
  2371 => x"921480f5",
  2372 => x"2d737081",
  2373 => x"055581b7",
  2374 => x"2d941480",
  2375 => x"f52d7370",
  2376 => x"81055581",
  2377 => x"b72d9614",
  2378 => x"80f52d73",
  2379 => x"70810555",
  2380 => x"81b72d98",
  2381 => x"1480f52d",
  2382 => x"73708105",
  2383 => x"5581b72d",
  2384 => x"9c1480f5",
  2385 => x"2d737081",
  2386 => x"055581b7",
  2387 => x"2d9e1480",
  2388 => x"f52d7381",
  2389 => x"b72d7780",
  2390 => x"da940c80",
  2391 => x"537280db",
  2392 => x"d00c02a0",
  2393 => x"050d0402",
  2394 => x"cc050d7e",
  2395 => x"605e5a80",
  2396 => x"0b80e3f8",
  2397 => x"0880e3fc",
  2398 => x"08595c56",
  2399 => x"805880e3",
  2400 => x"d808782e",
  2401 => x"81bc3877",
  2402 => x"8f06a017",
  2403 => x"57547391",
  2404 => x"3880ddc8",
  2405 => x"52765181",
  2406 => x"1757be85",
  2407 => x"2d80ddc8",
  2408 => x"56807680",
  2409 => x"f52d5654",
  2410 => x"74742e83",
  2411 => x"38815474",
  2412 => x"81e52e81",
  2413 => x"81388170",
  2414 => x"7506555c",
  2415 => x"73802e80",
  2416 => x"f5388b16",
  2417 => x"80f52d98",
  2418 => x"06597880",
  2419 => x"e9388b53",
  2420 => x"7c527551",
  2421 => x"bfa92d80",
  2422 => x"dbd00880",
  2423 => x"d9389c16",
  2424 => x"085180cd",
  2425 => x"e42d80db",
  2426 => x"d008841b",
  2427 => x"0c9a1680",
  2428 => x"e02d5180",
  2429 => x"ce952d80",
  2430 => x"dbd00880",
  2431 => x"dbd00888",
  2432 => x"1c0c80db",
  2433 => x"d0085555",
  2434 => x"80e3d408",
  2435 => x"802e9a38",
  2436 => x"941680e0",
  2437 => x"2d5180ce",
  2438 => x"952d80db",
  2439 => x"d008902b",
  2440 => x"83fff00a",
  2441 => x"06701651",
  2442 => x"5473881b",
  2443 => x"0c787a0c",
  2444 => x"7b5480cd",
  2445 => x"80048118",
  2446 => x"5880e3d8",
  2447 => x"087826fe",
  2448 => x"c63880e3",
  2449 => x"d408802e",
  2450 => x"b5387a51",
  2451 => x"80c7af2d",
  2452 => x"80dbd008",
  2453 => x"80dbd008",
  2454 => x"80ffffff",
  2455 => x"f806555b",
  2456 => x"7380ffff",
  2457 => x"fff82e96",
  2458 => x"3880dbd0",
  2459 => x"08fe0580",
  2460 => x"e3cc0829",
  2461 => x"80e3e008",
  2462 => x"055780ca",
  2463 => x"fc048054",
  2464 => x"7380dbd0",
  2465 => x"0c02b405",
  2466 => x"0d0402f4",
  2467 => x"050d7470",
  2468 => x"08810571",
  2469 => x"0c700880",
  2470 => x"e3d00806",
  2471 => x"53537190",
  2472 => x"38881308",
  2473 => x"5180c7af",
  2474 => x"2d80dbd0",
  2475 => x"0888140c",
  2476 => x"810b80db",
  2477 => x"d00c028c",
  2478 => x"050d0402",
  2479 => x"f0050d75",
  2480 => x"881108fe",
  2481 => x"0580e3cc",
  2482 => x"082980e3",
  2483 => x"e0081172",
  2484 => x"0880e3d0",
  2485 => x"08060579",
  2486 => x"55535454",
  2487 => x"be852d02",
  2488 => x"90050d04",
  2489 => x"02f4050d",
  2490 => x"7470882a",
  2491 => x"83fe8006",
  2492 => x"7072982a",
  2493 => x"0772882b",
  2494 => x"87fc8080",
  2495 => x"0673982b",
  2496 => x"81f00a06",
  2497 => x"71730707",
  2498 => x"80dbd00c",
  2499 => x"56515351",
  2500 => x"028c050d",
  2501 => x"0402f805",
  2502 => x"0d028e05",
  2503 => x"80f52d74",
  2504 => x"882b0770",
  2505 => x"83ffff06",
  2506 => x"80dbd00c",
  2507 => x"51028805",
  2508 => x"0d0402f4",
  2509 => x"050d7476",
  2510 => x"78535452",
  2511 => x"80712597",
  2512 => x"38727081",
  2513 => x"055480f5",
  2514 => x"2d727081",
  2515 => x"055481b7",
  2516 => x"2dff1151",
  2517 => x"70eb3880",
  2518 => x"7281b72d",
  2519 => x"028c050d",
  2520 => x"0402e805",
  2521 => x"0d775680",
  2522 => x"70565473",
  2523 => x"7624b738",
  2524 => x"80e3d808",
  2525 => x"742eaf38",
  2526 => x"735180c8",
  2527 => x"ab2d80db",
  2528 => x"d00880db",
  2529 => x"d0080981",
  2530 => x"057080db",
  2531 => x"d008079f",
  2532 => x"2a770581",
  2533 => x"17575753",
  2534 => x"53747624",
  2535 => x"893880e3",
  2536 => x"d8087426",
  2537 => x"d3387280",
  2538 => x"dbd00c02",
  2539 => x"98050d04",
  2540 => x"02f0050d",
  2541 => x"80dbcc08",
  2542 => x"165180ce",
  2543 => x"e12d80db",
  2544 => x"d008802e",
  2545 => x"a0388b53",
  2546 => x"80dbd008",
  2547 => x"5280e1c8",
  2548 => x"5180ceb2",
  2549 => x"2d80e484",
  2550 => x"08547380",
  2551 => x"2e873880",
  2552 => x"e1c85173",
  2553 => x"2d029005",
  2554 => x"0d0402dc",
  2555 => x"050d8070",
  2556 => x"5a557480",
  2557 => x"dbcc0825",
  2558 => x"b53880e3",
  2559 => x"d808752e",
  2560 => x"ad387851",
  2561 => x"80c8ab2d",
  2562 => x"80dbd008",
  2563 => x"09810570",
  2564 => x"80dbd008",
  2565 => x"079f2a76",
  2566 => x"05811b5b",
  2567 => x"56547480",
  2568 => x"dbcc0825",
  2569 => x"893880e3",
  2570 => x"d8087926",
  2571 => x"d5388055",
  2572 => x"7880e3d8",
  2573 => x"082781e4",
  2574 => x"38785180",
  2575 => x"c8ab2d80",
  2576 => x"dbd00880",
  2577 => x"2e81b438",
  2578 => x"80dbd008",
  2579 => x"8b0580f5",
  2580 => x"2d70842a",
  2581 => x"70810677",
  2582 => x"1078842b",
  2583 => x"80e1c80b",
  2584 => x"80f52d5c",
  2585 => x"5c535155",
  2586 => x"5673802e",
  2587 => x"80ce3874",
  2588 => x"16822b80",
  2589 => x"d2c00b80",
  2590 => x"daa0120c",
  2591 => x"54777531",
  2592 => x"1080e488",
  2593 => x"11555690",
  2594 => x"74708105",
  2595 => x"5681b72d",
  2596 => x"a07481b7",
  2597 => x"2d7681ff",
  2598 => x"06811658",
  2599 => x"5473802e",
  2600 => x"8b389c53",
  2601 => x"80e1c852",
  2602 => x"80d1b304",
  2603 => x"8b5380db",
  2604 => x"d0085280",
  2605 => x"e48a1651",
  2606 => x"80d1f104",
  2607 => x"7416822b",
  2608 => x"80cfb00b",
  2609 => x"80daa012",
  2610 => x"0c547681",
  2611 => x"ff068116",
  2612 => x"58547380",
  2613 => x"2e8b389c",
  2614 => x"5380e1c8",
  2615 => x"5280d1e8",
  2616 => x"048b5380",
  2617 => x"dbd00852",
  2618 => x"77753110",
  2619 => x"80e48805",
  2620 => x"51765580",
  2621 => x"ceb22d80",
  2622 => x"d2900474",
  2623 => x"90297531",
  2624 => x"701080e4",
  2625 => x"88055154",
  2626 => x"80dbd008",
  2627 => x"7481b72d",
  2628 => x"81195974",
  2629 => x"8b24a438",
  2630 => x"80d0b004",
  2631 => x"74902975",
  2632 => x"31701080",
  2633 => x"e488058c",
  2634 => x"77315751",
  2635 => x"54807481",
  2636 => x"b72d9e14",
  2637 => x"ff165654",
  2638 => x"74f33802",
  2639 => x"a4050d04",
  2640 => x"02fc050d",
  2641 => x"80dbcc08",
  2642 => x"135180ce",
  2643 => x"e12d80db",
  2644 => x"d008802e",
  2645 => x"893880db",
  2646 => x"d00851bf",
  2647 => x"e82d800b",
  2648 => x"80dbcc0c",
  2649 => x"80cfea2d",
  2650 => x"adf22d02",
  2651 => x"84050d04",
  2652 => x"02fc050d",
  2653 => x"725170fd",
  2654 => x"2eb23870",
  2655 => x"fd248b38",
  2656 => x"70fc2e80",
  2657 => x"d03880d3",
  2658 => x"df0470fe",
  2659 => x"2eb93870",
  2660 => x"ff2e0981",
  2661 => x"0680c838",
  2662 => x"80dbcc08",
  2663 => x"5170802e",
  2664 => x"be38ff11",
  2665 => x"80dbcc0c",
  2666 => x"80d3df04",
  2667 => x"80dbcc08",
  2668 => x"f0057080",
  2669 => x"dbcc0c51",
  2670 => x"708025a3",
  2671 => x"38800b80",
  2672 => x"dbcc0c80",
  2673 => x"d3df0480",
  2674 => x"dbcc0881",
  2675 => x"0580dbcc",
  2676 => x"0c80d3df",
  2677 => x"0480dbcc",
  2678 => x"08900580",
  2679 => x"dbcc0c80",
  2680 => x"cfea2dad",
  2681 => x"f22d0284",
  2682 => x"050d0402",
  2683 => x"fc050d80",
  2684 => x"0b80dbcc",
  2685 => x"0c80cfea",
  2686 => x"2dacee2d",
  2687 => x"80dbd008",
  2688 => x"80dbbc0c",
  2689 => x"80da9851",
  2690 => x"af982d02",
  2691 => x"84050d04",
  2692 => x"7180e484",
  2693 => x"0c040000",
  2694 => x"00ffffff",
  2695 => x"ff00ffff",
  2696 => x"ffff00ff",
  2697 => x"ffffff00",
  2698 => x"30313233",
  2699 => x"34353637",
  2700 => x"38394142",
  2701 => x"43444546",
  2702 => x"00000000",
  2703 => x"44656275",
  2704 => x"67000000",
  2705 => x"52657365",
  2706 => x"74000000",
  2707 => x"5363616e",
  2708 => x"6c696e65",
  2709 => x"73000000",
  2710 => x"50414c20",
  2711 => x"2f204e54",
  2712 => x"53430000",
  2713 => x"436f6c6f",
  2714 => x"72000000",
  2715 => x"44696666",
  2716 => x"6963756c",
  2717 => x"74792041",
  2718 => x"00000000",
  2719 => x"44696666",
  2720 => x"6963756c",
  2721 => x"74792042",
  2722 => x"00000000",
  2723 => x"53757065",
  2724 => x"72636869",
  2725 => x"7020696e",
  2726 => x"20636172",
  2727 => x"74726964",
  2728 => x"67650000",
  2729 => x"524f4d00",
  2730 => x"626f6f74",
  2731 => x"00000000",
  2732 => x"53656c65",
  2733 => x"63740000",
  2734 => x"53746172",
  2735 => x"74000000",
  2736 => x"4c6f6164",
  2737 => x"20524f4d",
  2738 => x"20100000",
  2739 => x"45786974",
  2740 => x"00000000",
  2741 => x"524f4d20",
  2742 => x"6c6f6164",
  2743 => x"696e6720",
  2744 => x"6661696c",
  2745 => x"65640000",
  2746 => x"4f4b0000",
  2747 => x"45525220",
  2748 => x"00000000",
  2749 => x"496e6974",
  2750 => x"69616c69",
  2751 => x"7a696e67",
  2752 => x"20534420",
  2753 => x"63617264",
  2754 => x"0a000000",
  2755 => x"436f6c6c",
  2756 => x"6563746f",
  2757 => x"72566973",
  2758 => x"696f6e00",
  2759 => x"16200000",
  2760 => x"14200000",
  2761 => x"15200000",
  2762 => x"53442069",
  2763 => x"6e69742e",
  2764 => x"2e2e0a00",
  2765 => x"53442063",
  2766 => x"61726420",
  2767 => x"72657365",
  2768 => x"74206661",
  2769 => x"696c6564",
  2770 => x"210a0000",
  2771 => x"53444843",
  2772 => x"20657272",
  2773 => x"6f72210a",
  2774 => x"00000000",
  2775 => x"57726974",
  2776 => x"65206661",
  2777 => x"696c6564",
  2778 => x"0a000000",
  2779 => x"52656164",
  2780 => x"20666169",
  2781 => x"6c65640a",
  2782 => x"00000000",
  2783 => x"43617264",
  2784 => x"20696e69",
  2785 => x"74206661",
  2786 => x"696c6564",
  2787 => x"0a000000",
  2788 => x"46415431",
  2789 => x"36202020",
  2790 => x"00000000",
  2791 => x"46415433",
  2792 => x"32202020",
  2793 => x"00000000",
  2794 => x"4e6f2070",
  2795 => x"61727469",
  2796 => x"74696f6e",
  2797 => x"20736967",
  2798 => x"0a000000",
  2799 => x"42616420",
  2800 => x"70617274",
  2801 => x"0a000000",
  2802 => x"4261636b",
  2803 => x"00000000",
  2804 => x"00000002",
  2805 => x"00002a28",
  2806 => x"00002e3c",
  2807 => x"00000002",
  2808 => x"00002df8",
  2809 => x"0000138d",
  2810 => x"00000002",
  2811 => x"00002a3c",
  2812 => x"00001321",
  2813 => x"00000002",
  2814 => x"00002a44",
  2815 => x"0000035a",
  2816 => x"00000001",
  2817 => x"00002a4c",
  2818 => x"00000000",
  2819 => x"00000001",
  2820 => x"00002a58",
  2821 => x"00000001",
  2822 => x"00000001",
  2823 => x"00002a64",
  2824 => x"00000002",
  2825 => x"00000001",
  2826 => x"00002a6c",
  2827 => x"00000003",
  2828 => x"00000001",
  2829 => x"00002a7c",
  2830 => x"00000004",
  2831 => x"00000001",
  2832 => x"00002a8c",
  2833 => x"00000005",
  2834 => x"00000001",
  2835 => x"00002aa4",
  2836 => x"00000006",
  2837 => x"00000002",
  2838 => x"00002aa8",
  2839 => x"00001110",
  2840 => x"00000002",
  2841 => x"00002ab0",
  2842 => x"0000036e",
  2843 => x"00000002",
  2844 => x"00002ab8",
  2845 => x"00000a3f",
  2846 => x"00000002",
  2847 => x"00002ac0",
  2848 => x"000029eb",
  2849 => x"00000002",
  2850 => x"00002acc",
  2851 => x"0000168b",
  2852 => x"00000000",
  2853 => x"00000000",
  2854 => x"00000000",
  2855 => x"00000004",
  2856 => x"00002ad4",
  2857 => x"00002c9c",
  2858 => x"00000004",
  2859 => x"00002ae8",
  2860 => x"00002bdc",
  2861 => x"00000000",
  2862 => x"00000000",
  2863 => x"00000000",
  2864 => x"00000000",
  2865 => x"00000000",
  2866 => x"00000000",
  2867 => x"00000000",
  2868 => x"00000000",
  2869 => x"00000000",
  2870 => x"00000000",
  2871 => x"00000000",
  2872 => x"00000000",
  2873 => x"00000000",
  2874 => x"00000000",
  2875 => x"00000000",
  2876 => x"00000000",
  2877 => x"00000000",
  2878 => x"00000000",
  2879 => x"00000000",
  2880 => x"00000000",
  2881 => x"00000000",
  2882 => x"00000000",
  2883 => x"00000006",
  2884 => x"00000000",
  2885 => x"00000000",
  2886 => x"00000002",
  2887 => x"00003208",
  2888 => x"000027b0",
  2889 => x"00000002",
  2890 => x"00003226",
  2891 => x"000027b0",
  2892 => x"00000002",
  2893 => x"00003244",
  2894 => x"000027b0",
  2895 => x"00000002",
  2896 => x"00003262",
  2897 => x"000027b0",
  2898 => x"00000002",
  2899 => x"00003280",
  2900 => x"000027b0",
  2901 => x"00000002",
  2902 => x"0000329e",
  2903 => x"000027b0",
  2904 => x"00000002",
  2905 => x"000032bc",
  2906 => x"000027b0",
  2907 => x"00000002",
  2908 => x"000032da",
  2909 => x"000027b0",
  2910 => x"00000002",
  2911 => x"000032f8",
  2912 => x"000027b0",
  2913 => x"00000002",
  2914 => x"00003316",
  2915 => x"000027b0",
  2916 => x"00000002",
  2917 => x"00003334",
  2918 => x"000027b0",
  2919 => x"00000002",
  2920 => x"00003352",
  2921 => x"000027b0",
  2922 => x"00000002",
  2923 => x"00003370",
  2924 => x"000027b0",
  2925 => x"00000004",
  2926 => x"00002bc8",
  2927 => x"00000000",
  2928 => x"00000000",
  2929 => x"00000000",
  2930 => x"00002970",
  2931 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

