-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80e2",
     9 => x"9c080b0b",
    10 => x"80e2a008",
    11 => x"0b0b80e2",
    12 => x"a4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"e2a40c0b",
    16 => x"0b80e2a0",
    17 => x"0c0b0b80",
    18 => x"e29c0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d9bc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80e29c70",
    57 => x"80edd427",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a797",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80e2",
    65 => x"ac0c9f0b",
    66 => x"80e2b00c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"e2b008ff",
    70 => x"0580e2b0",
    71 => x"0c80e2b0",
    72 => x"088025e8",
    73 => x"3880e2ac",
    74 => x"08ff0580",
    75 => x"e2ac0c80",
    76 => x"e2ac0880",
    77 => x"25d03880",
    78 => x"0b80e2b0",
    79 => x"0c800b80",
    80 => x"e2ac0c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80e2ac08",
   100 => x"25913882",
   101 => x"c82d80e2",
   102 => x"ac08ff05",
   103 => x"80e2ac0c",
   104 => x"838a0480",
   105 => x"e2ac0880",
   106 => x"e2b00853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80e2ac08",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"e2b00881",
   116 => x"0580e2b0",
   117 => x"0c80e2b0",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80e2b0",
   121 => x"0c80e2ac",
   122 => x"08810580",
   123 => x"e2ac0c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480e2",
   128 => x"b0088105",
   129 => x"80e2b00c",
   130 => x"80e2b008",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80e2b0",
   134 => x"0c80e2ac",
   135 => x"08810580",
   136 => x"e2ac0c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"e2b40cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"e2b40c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280e2",
   177 => x"b4088407",
   178 => x"80e2b40c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80dd",
   183 => x"9c0c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80e2b4",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80e2",
   208 => x"9c0c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02fc050d",
  1093 => x"ffb40870",
  1094 => x"9f2a80e2",
  1095 => x"9c0c5102",
  1096 => x"84050d04",
  1097 => x"02f4050d",
  1098 => x"a2902d80",
  1099 => x"e0ac0886",
  1100 => x"2a80e29c",
  1101 => x"08822b84",
  1102 => x"32718106",
  1103 => x"07708207",
  1104 => x"e00c5152",
  1105 => x"805186da",
  1106 => x"2d028c05",
  1107 => x"0d0402f4",
  1108 => x"050d7476",
  1109 => x"54527270",
  1110 => x"81055480",
  1111 => x"f52d5170",
  1112 => x"72708105",
  1113 => x"5481b72d",
  1114 => x"70ec3870",
  1115 => x"7281b72d",
  1116 => x"028c050d",
  1117 => x"0402f405",
  1118 => x"0d80ddb8",
  1119 => x"0b80f52d",
  1120 => x"80e0ac08",
  1121 => x"70810653",
  1122 => x"54527080",
  1123 => x"2e853871",
  1124 => x"84075272",
  1125 => x"812a7081",
  1126 => x"06515170",
  1127 => x"802e8538",
  1128 => x"71820752",
  1129 => x"72822a70",
  1130 => x"81065151",
  1131 => x"70802e85",
  1132 => x"38718107",
  1133 => x"5272832a",
  1134 => x"70810651",
  1135 => x"5170802e",
  1136 => x"85387188",
  1137 => x"07527284",
  1138 => x"2a708106",
  1139 => x"51517080",
  1140 => x"2e853871",
  1141 => x"90075272",
  1142 => x"852a7081",
  1143 => x"06515170",
  1144 => x"802e8538",
  1145 => x"71a00752",
  1146 => x"72882a70",
  1147 => x"81065151",
  1148 => x"70802e86",
  1149 => x"387180c0",
  1150 => x"07527289",
  1151 => x"2a708106",
  1152 => x"51517080",
  1153 => x"2e863871",
  1154 => x"81800752",
  1155 => x"71fc0c71",
  1156 => x"80e29c0c",
  1157 => x"028c050d",
  1158 => x"0402cc05",
  1159 => x"0d7e5d80",
  1160 => x"0b80e0ac",
  1161 => x"08818006",
  1162 => x"715c5d5b",
  1163 => x"810bec0c",
  1164 => x"840bec0c",
  1165 => x"7c5280e2",
  1166 => x"b85180ce",
  1167 => x"df2d80e2",
  1168 => x"9c087b2e",
  1169 => x"80ff3880",
  1170 => x"e2bc087b",
  1171 => x"ff125759",
  1172 => x"57747b2e",
  1173 => x"8b388118",
  1174 => x"75812a56",
  1175 => x"5874f738",
  1176 => x"f7185881",
  1177 => x"5b807725",
  1178 => x"80db3877",
  1179 => x"52745184",
  1180 => x"a82d80e3",
  1181 => x"8c5280e2",
  1182 => x"b85180d1",
  1183 => x"b52d80e2",
  1184 => x"9c08802e",
  1185 => x"a63880e3",
  1186 => x"8c597ba7",
  1187 => x"3883ff56",
  1188 => x"78708105",
  1189 => x"5a80f52d",
  1190 => x"7a811c5c",
  1191 => x"e40ce80c",
  1192 => x"ff165675",
  1193 => x"8025e938",
  1194 => x"a5b30480",
  1195 => x"e29c085b",
  1196 => x"84805780",
  1197 => x"e2b85180",
  1198 => x"d1842dfc",
  1199 => x"80178116",
  1200 => x"5657a4e5",
  1201 => x"0480e2bc",
  1202 => x"08f80c88",
  1203 => x"1d548074",
  1204 => x"80f52d70",
  1205 => x"81ff0655",
  1206 => x"58557275",
  1207 => x"2eb63881",
  1208 => x"1480f52d",
  1209 => x"5372752e",
  1210 => x"ab387482",
  1211 => x"1580f52d",
  1212 => x"54567280",
  1213 => x"d32e0981",
  1214 => x"06833881",
  1215 => x"567280f3",
  1216 => x"32700981",
  1217 => x"05708025",
  1218 => x"78075151",
  1219 => x"5372802e",
  1220 => x"8338a055",
  1221 => x"807781ff",
  1222 => x"06545672",
  1223 => x"80c52e09",
  1224 => x"81068338",
  1225 => x"81567280",
  1226 => x"e5327009",
  1227 => x"81057080",
  1228 => x"25780751",
  1229 => x"51537280",
  1230 => x"2ea43881",
  1231 => x"1480f52d",
  1232 => x"5372b02e",
  1233 => x"09810689",
  1234 => x"38748280",
  1235 => x"0755a6de",
  1236 => x"0472b72e",
  1237 => x"09810686",
  1238 => x"38748480",
  1239 => x"075580e0",
  1240 => x"ac08f9df",
  1241 => x"06750780",
  1242 => x"e0ac0ca2",
  1243 => x"f52d800b",
  1244 => x"e00c8051",
  1245 => x"86da2d86",
  1246 => x"c72d7a80",
  1247 => x"2e883880",
  1248 => x"dda451a7",
  1249 => x"8a0480de",
  1250 => x"d851b1a3",
  1251 => x"2d7a80e2",
  1252 => x"9c0c02b4",
  1253 => x"050d0402",
  1254 => x"f4050d84",
  1255 => x"0bec0ca2",
  1256 => x"902d80e2",
  1257 => x"9c08822b",
  1258 => x"8107e00c",
  1259 => x"aee02da8",
  1260 => x"ba2d81f9",
  1261 => x"2d8352ae",
  1262 => x"c32d8151",
  1263 => x"858d2dff",
  1264 => x"12527180",
  1265 => x"25f13884",
  1266 => x"0bec0c80",
  1267 => x"dba05186",
  1268 => x"a02d80c3",
  1269 => x"b72d80e2",
  1270 => x"9c08802e",
  1271 => x"80c53880",
  1272 => x"dbb85186",
  1273 => x"a02da499",
  1274 => x"5180d9b6",
  1275 => x"2d80dda4",
  1276 => x"51b1a32d",
  1277 => x"af822da9",
  1278 => x"e52d80e2",
  1279 => x"9c088106",
  1280 => x"5271802e",
  1281 => x"86388051",
  1282 => x"94bf2db1",
  1283 => x"b62d80e2",
  1284 => x"9c0852a2",
  1285 => x"f52d8653",
  1286 => x"71833884",
  1287 => x"5372ec0c",
  1288 => x"a7f70480",
  1289 => x"0b80e29c",
  1290 => x"0c028c05",
  1291 => x"0d047198",
  1292 => x"0c04ffb0",
  1293 => x"0880e29c",
  1294 => x"0c04810b",
  1295 => x"ffb00c04",
  1296 => x"800bffb0",
  1297 => x"0c0402d8",
  1298 => x"050dffb4",
  1299 => x"0887ffff",
  1300 => x"065a8154",
  1301 => x"807080e0",
  1302 => x"980880e0",
  1303 => x"9c0880df",
  1304 => x"f45b5957",
  1305 => x"5a587974",
  1306 => x"06757506",
  1307 => x"52527171",
  1308 => x"2e8d3880",
  1309 => x"77818a2d",
  1310 => x"73097506",
  1311 => x"72075576",
  1312 => x"80e02d70",
  1313 => x"83ffff06",
  1314 => x"53517180",
  1315 => x"e42e0981",
  1316 => x"06a23874",
  1317 => x"74067077",
  1318 => x"76063270",
  1319 => x"09810570",
  1320 => x"72079f2a",
  1321 => x"7b057709",
  1322 => x"7a067407",
  1323 => x"5a5b5353",
  1324 => x"53a9c204",
  1325 => x"7180e426",
  1326 => x"89388111",
  1327 => x"51707781",
  1328 => x"8a2d7310",
  1329 => x"811a8219",
  1330 => x"595a5490",
  1331 => x"7925ff96",
  1332 => x"387580e0",
  1333 => x"9c0c7480",
  1334 => x"e0980c77",
  1335 => x"80e29c0c",
  1336 => x"02a8050d",
  1337 => x"0402d005",
  1338 => x"0d805caa",
  1339 => x"f50480e2",
  1340 => x"9c0881f0",
  1341 => x"2e098106",
  1342 => x"8a38810b",
  1343 => x"80e0a40c",
  1344 => x"aaf50480",
  1345 => x"e29c0881",
  1346 => x"e02e0981",
  1347 => x"068a3881",
  1348 => x"0b80e0a8",
  1349 => x"0caaf504",
  1350 => x"80e29c08",
  1351 => x"5280e0a8",
  1352 => x"08802e89",
  1353 => x"3880e29c",
  1354 => x"08818005",
  1355 => x"5271842c",
  1356 => x"728f0653",
  1357 => x"5380e0a4",
  1358 => x"08802e9a",
  1359 => x"38728429",
  1360 => x"80defc05",
  1361 => x"72138171",
  1362 => x"2b700973",
  1363 => x"0806730c",
  1364 => x"515353aa",
  1365 => x"e9047284",
  1366 => x"2980defc",
  1367 => x"05721383",
  1368 => x"712b7208",
  1369 => x"07720c53",
  1370 => x"53800b80",
  1371 => x"e0a80c80",
  1372 => x"0b80e0a4",
  1373 => x"0c80e2c4",
  1374 => x"51adb62d",
  1375 => x"80e29c08",
  1376 => x"ff24feea",
  1377 => x"38a8c62d",
  1378 => x"80e29c08",
  1379 => x"802e81b0",
  1380 => x"38815980",
  1381 => x"0b80e0a0",
  1382 => x"0880e09c",
  1383 => x"0880dfd0",
  1384 => x"5a5c5c58",
  1385 => x"7a79067a",
  1386 => x"7a065452",
  1387 => x"71732e80",
  1388 => x"f8387209",
  1389 => x"81057074",
  1390 => x"07802580",
  1391 => x"dfbc1a80",
  1392 => x"f52d7084",
  1393 => x"2c718f06",
  1394 => x"58535757",
  1395 => x"5275802e",
  1396 => x"a3387184",
  1397 => x"2980defc",
  1398 => x"05741583",
  1399 => x"712b7208",
  1400 => x"07720c54",
  1401 => x"527680e0",
  1402 => x"2d810552",
  1403 => x"7177818a",
  1404 => x"2dac8a04",
  1405 => x"71842980",
  1406 => x"defc0574",
  1407 => x"1581712b",
  1408 => x"70097308",
  1409 => x"06730c51",
  1410 => x"53537485",
  1411 => x"32700981",
  1412 => x"05708025",
  1413 => x"51515275",
  1414 => x"802e8e38",
  1415 => x"81707306",
  1416 => x"53537180",
  1417 => x"2e833872",
  1418 => x"5c781081",
  1419 => x"19821959",
  1420 => x"59599078",
  1421 => x"25feed38",
  1422 => x"80e09c08",
  1423 => x"80e0a00c",
  1424 => x"7b80e29c",
  1425 => x"0c02b005",
  1426 => x"0d0402f8",
  1427 => x"050d80de",
  1428 => x"fc528f51",
  1429 => x"80727084",
  1430 => x"05540cff",
  1431 => x"11517080",
  1432 => x"25f23802",
  1433 => x"88050d04",
  1434 => x"02f0050d",
  1435 => x"7551a8c0",
  1436 => x"2d70822c",
  1437 => x"fc0680de",
  1438 => x"fc117210",
  1439 => x"9e067108",
  1440 => x"70722a70",
  1441 => x"83068274",
  1442 => x"2b700974",
  1443 => x"06760c54",
  1444 => x"51565753",
  1445 => x"5153a8ba",
  1446 => x"2d7180e2",
  1447 => x"9c0c0290",
  1448 => x"050d0402",
  1449 => x"fc050d72",
  1450 => x"5180710c",
  1451 => x"800b8412",
  1452 => x"0c028405",
  1453 => x"0d0402f0",
  1454 => x"050d7570",
  1455 => x"08841208",
  1456 => x"535353ff",
  1457 => x"5471712e",
  1458 => x"a838a8c0",
  1459 => x"2d841308",
  1460 => x"70842914",
  1461 => x"88117008",
  1462 => x"7081ff06",
  1463 => x"84180881",
  1464 => x"11870684",
  1465 => x"1a0c5351",
  1466 => x"55515151",
  1467 => x"a8ba2d71",
  1468 => x"547380e2",
  1469 => x"9c0c0290",
  1470 => x"050d0402",
  1471 => x"f8050da8",
  1472 => x"c02de008",
  1473 => x"708b2a70",
  1474 => x"81065152",
  1475 => x"5270802e",
  1476 => x"a13880e2",
  1477 => x"c4087084",
  1478 => x"2980e2cc",
  1479 => x"057381ff",
  1480 => x"06710c51",
  1481 => x"5180e2c4",
  1482 => x"08811187",
  1483 => x"0680e2c4",
  1484 => x"0c51800b",
  1485 => x"80e2ec0c",
  1486 => x"a8b22da8",
  1487 => x"ba2d0288",
  1488 => x"050d0402",
  1489 => x"fc050da8",
  1490 => x"c02d810b",
  1491 => x"80e2ec0c",
  1492 => x"a8ba2d80",
  1493 => x"e2ec0851",
  1494 => x"70f93802",
  1495 => x"84050d04",
  1496 => x"02fc050d",
  1497 => x"80e2c451",
  1498 => x"ada32dac",
  1499 => x"ca2dadfb",
  1500 => x"51a8ae2d",
  1501 => x"0284050d",
  1502 => x"0480e2f8",
  1503 => x"0880e29c",
  1504 => x"0c0402fc",
  1505 => x"050d810b",
  1506 => x"80e0b00c",
  1507 => x"8151858d",
  1508 => x"2d028405",
  1509 => x"0d0402fc",
  1510 => x"050dafa0",
  1511 => x"04a9e52d",
  1512 => x"80f651ac",
  1513 => x"e82d80e2",
  1514 => x"9c08f238",
  1515 => x"80da51ac",
  1516 => x"e82d80e2",
  1517 => x"9c08e638",
  1518 => x"80e29c08",
  1519 => x"80e0b00c",
  1520 => x"80e29c08",
  1521 => x"51858d2d",
  1522 => x"0284050d",
  1523 => x"0402ec05",
  1524 => x"0d765480",
  1525 => x"52870b88",
  1526 => x"1580f52d",
  1527 => x"56537472",
  1528 => x"248338a0",
  1529 => x"53725183",
  1530 => x"842d8112",
  1531 => x"8b1580f5",
  1532 => x"2d545272",
  1533 => x"7225de38",
  1534 => x"0294050d",
  1535 => x"0402f005",
  1536 => x"0d80e2f8",
  1537 => x"085481f9",
  1538 => x"2d800b80",
  1539 => x"e2fc0c73",
  1540 => x"08802e81",
  1541 => x"8938820b",
  1542 => x"80e2b00c",
  1543 => x"80e2fc08",
  1544 => x"8f0680e2",
  1545 => x"ac0c7308",
  1546 => x"5271832e",
  1547 => x"96387183",
  1548 => x"26893871",
  1549 => x"812eb038",
  1550 => x"b1870471",
  1551 => x"852ea038",
  1552 => x"b1870488",
  1553 => x"1480f52d",
  1554 => x"84150880",
  1555 => x"dbd05354",
  1556 => x"5286a02d",
  1557 => x"71842913",
  1558 => x"70085252",
  1559 => x"b18b0473",
  1560 => x"51afcd2d",
  1561 => x"b1870480",
  1562 => x"e0ac0888",
  1563 => x"15082c70",
  1564 => x"81065152",
  1565 => x"71802e88",
  1566 => x"3880dbd4",
  1567 => x"51b18404",
  1568 => x"80dbd851",
  1569 => x"86a02d84",
  1570 => x"14085186",
  1571 => x"a02d80e2",
  1572 => x"fc088105",
  1573 => x"80e2fc0c",
  1574 => x"8c1454b0",
  1575 => x"8f040290",
  1576 => x"050d0471",
  1577 => x"80e2f80c",
  1578 => x"affd2d80",
  1579 => x"e2fc08ff",
  1580 => x"0580e380",
  1581 => x"0c0402e8",
  1582 => x"050d80e2",
  1583 => x"f80880e3",
  1584 => x"84085755",
  1585 => x"80f651ac",
  1586 => x"e82d80e2",
  1587 => x"9c08812a",
  1588 => x"70810651",
  1589 => x"5271802e",
  1590 => x"a438b1e0",
  1591 => x"04a9e52d",
  1592 => x"80f651ac",
  1593 => x"e82d80e2",
  1594 => x"9c08f238",
  1595 => x"80e0b008",
  1596 => x"81327080",
  1597 => x"e0b00c70",
  1598 => x"5252858d",
  1599 => x"2d800b80",
  1600 => x"e2f00c80",
  1601 => x"0b80e2f4",
  1602 => x"0c80e0b0",
  1603 => x"08838d38",
  1604 => x"80da51ac",
  1605 => x"e82d80e2",
  1606 => x"9c08802e",
  1607 => x"8c3880e2",
  1608 => x"f0088180",
  1609 => x"0780e2f0",
  1610 => x"0c80d951",
  1611 => x"ace82d80",
  1612 => x"e29c0880",
  1613 => x"2e8c3880",
  1614 => x"e2f00880",
  1615 => x"c00780e2",
  1616 => x"f00c8194",
  1617 => x"51ace82d",
  1618 => x"80e29c08",
  1619 => x"802e8b38",
  1620 => x"80e2f008",
  1621 => x"900780e2",
  1622 => x"f00c8191",
  1623 => x"51ace82d",
  1624 => x"80e29c08",
  1625 => x"802e8b38",
  1626 => x"80e2f008",
  1627 => x"a00780e2",
  1628 => x"f00c81f5",
  1629 => x"51ace82d",
  1630 => x"80e29c08",
  1631 => x"802e8b38",
  1632 => x"80e2f008",
  1633 => x"810780e2",
  1634 => x"f00c81f2",
  1635 => x"51ace82d",
  1636 => x"80e29c08",
  1637 => x"802e8b38",
  1638 => x"80e2f008",
  1639 => x"820780e2",
  1640 => x"f00c81eb",
  1641 => x"51ace82d",
  1642 => x"80e29c08",
  1643 => x"802e8b38",
  1644 => x"80e2f008",
  1645 => x"840780e2",
  1646 => x"f00c81f4",
  1647 => x"51ace82d",
  1648 => x"80e29c08",
  1649 => x"802e8b38",
  1650 => x"80e2f008",
  1651 => x"880780e2",
  1652 => x"f00c80d8",
  1653 => x"51ace82d",
  1654 => x"80e29c08",
  1655 => x"802e8c38",
  1656 => x"80e2f408",
  1657 => x"81800780",
  1658 => x"e2f40c92",
  1659 => x"51ace82d",
  1660 => x"80e29c08",
  1661 => x"802e8c38",
  1662 => x"80e2f408",
  1663 => x"80c00780",
  1664 => x"e2f40c94",
  1665 => x"51ace82d",
  1666 => x"80e29c08",
  1667 => x"802e8b38",
  1668 => x"80e2f408",
  1669 => x"900780e2",
  1670 => x"f40c9151",
  1671 => x"ace82d80",
  1672 => x"e29c0880",
  1673 => x"2e8b3880",
  1674 => x"e2f408a0",
  1675 => x"0780e2f4",
  1676 => x"0c9d51ac",
  1677 => x"e82d80e2",
  1678 => x"9c08802e",
  1679 => x"8b3880e2",
  1680 => x"f4088107",
  1681 => x"80e2f40c",
  1682 => x"9b51ace8",
  1683 => x"2d80e29c",
  1684 => x"08802e8b",
  1685 => x"3880e2f4",
  1686 => x"08820780",
  1687 => x"e2f40c9c",
  1688 => x"51ace82d",
  1689 => x"80e29c08",
  1690 => x"802e8b38",
  1691 => x"80e2f408",
  1692 => x"840780e2",
  1693 => x"f40ca351",
  1694 => x"ace82d80",
  1695 => x"e29c0880",
  1696 => x"2e8b3880",
  1697 => x"e2f40888",
  1698 => x"0780e2f4",
  1699 => x"0c81fd51",
  1700 => x"ace82d81",
  1701 => x"fa51ace8",
  1702 => x"2dbaf104",
  1703 => x"81f551ac",
  1704 => x"e82d80e2",
  1705 => x"9c08812a",
  1706 => x"70810651",
  1707 => x"5271802e",
  1708 => x"b33880e3",
  1709 => x"80085271",
  1710 => x"802e8a38",
  1711 => x"ff1280e3",
  1712 => x"800cb5e4",
  1713 => x"0480e2fc",
  1714 => x"081080e2",
  1715 => x"fc080570",
  1716 => x"84291651",
  1717 => x"52881208",
  1718 => x"802e8938",
  1719 => x"ff518812",
  1720 => x"0852712d",
  1721 => x"81f251ac",
  1722 => x"e82d80e2",
  1723 => x"9c08812a",
  1724 => x"70810651",
  1725 => x"5271802e",
  1726 => x"b43880e2",
  1727 => x"fc08ff11",
  1728 => x"80e38008",
  1729 => x"56535373",
  1730 => x"72258a38",
  1731 => x"811480e3",
  1732 => x"800cb6ad",
  1733 => x"04721013",
  1734 => x"70842916",
  1735 => x"51528812",
  1736 => x"08802e89",
  1737 => x"38fe5188",
  1738 => x"12085271",
  1739 => x"2d81fd51",
  1740 => x"ace82d80",
  1741 => x"e29c0881",
  1742 => x"2a708106",
  1743 => x"51527180",
  1744 => x"2eb13880",
  1745 => x"e3800880",
  1746 => x"2e8a3880",
  1747 => x"0b80e380",
  1748 => x"0cb6f304",
  1749 => x"80e2fc08",
  1750 => x"1080e2fc",
  1751 => x"08057084",
  1752 => x"29165152",
  1753 => x"88120880",
  1754 => x"2e8938fd",
  1755 => x"51881208",
  1756 => x"52712d81",
  1757 => x"fa51ace8",
  1758 => x"2d80e29c",
  1759 => x"08812a70",
  1760 => x"81065152",
  1761 => x"71802eb1",
  1762 => x"3880e2fc",
  1763 => x"08ff1154",
  1764 => x"5280e380",
  1765 => x"08732589",
  1766 => x"387280e3",
  1767 => x"800cb7b9",
  1768 => x"04711012",
  1769 => x"70842916",
  1770 => x"51528812",
  1771 => x"08802e89",
  1772 => x"38fc5188",
  1773 => x"12085271",
  1774 => x"2d80e380",
  1775 => x"08705354",
  1776 => x"73802e8a",
  1777 => x"388c15ff",
  1778 => x"155555b7",
  1779 => x"c004820b",
  1780 => x"80e2b00c",
  1781 => x"718f0680",
  1782 => x"e2ac0c81",
  1783 => x"eb51ace8",
  1784 => x"2d80e29c",
  1785 => x"08812a70",
  1786 => x"81065152",
  1787 => x"71802ead",
  1788 => x"38740885",
  1789 => x"2e098106",
  1790 => x"a4388815",
  1791 => x"80f52dff",
  1792 => x"05527188",
  1793 => x"1681b72d",
  1794 => x"71982b52",
  1795 => x"71802588",
  1796 => x"38800b88",
  1797 => x"1681b72d",
  1798 => x"7451afcd",
  1799 => x"2d81f451",
  1800 => x"ace82d80",
  1801 => x"e29c0881",
  1802 => x"2a708106",
  1803 => x"51527180",
  1804 => x"2eb33874",
  1805 => x"08852e09",
  1806 => x"8106aa38",
  1807 => x"881580f5",
  1808 => x"2d810552",
  1809 => x"71881681",
  1810 => x"b72d7181",
  1811 => x"ff068b16",
  1812 => x"80f52d54",
  1813 => x"52727227",
  1814 => x"87387288",
  1815 => x"1681b72d",
  1816 => x"7451afcd",
  1817 => x"2d80da51",
  1818 => x"ace82d80",
  1819 => x"e29c0881",
  1820 => x"2a708106",
  1821 => x"51527180",
  1822 => x"2e81ad38",
  1823 => x"80e2f808",
  1824 => x"80e38008",
  1825 => x"55537380",
  1826 => x"2e8a388c",
  1827 => x"13ff1555",
  1828 => x"53b98604",
  1829 => x"72085271",
  1830 => x"822ea638",
  1831 => x"71822689",
  1832 => x"3871812e",
  1833 => x"aa38baa8",
  1834 => x"0471832e",
  1835 => x"b4387184",
  1836 => x"2e098106",
  1837 => x"80f23888",
  1838 => x"130851b1",
  1839 => x"a32dbaa8",
  1840 => x"0480e380",
  1841 => x"08518813",
  1842 => x"0852712d",
  1843 => x"baa80481",
  1844 => x"0b881408",
  1845 => x"2b80e0ac",
  1846 => x"083280e0",
  1847 => x"ac0cb9fc",
  1848 => x"04881380",
  1849 => x"f52d8105",
  1850 => x"8b1480f5",
  1851 => x"2d535471",
  1852 => x"74248338",
  1853 => x"80547388",
  1854 => x"1481b72d",
  1855 => x"affd2dba",
  1856 => x"a8047508",
  1857 => x"802ea438",
  1858 => x"750851ac",
  1859 => x"e82d80e2",
  1860 => x"9c088106",
  1861 => x"5271802e",
  1862 => x"8c3880e3",
  1863 => x"80085184",
  1864 => x"16085271",
  1865 => x"2d881656",
  1866 => x"75d83880",
  1867 => x"54800b80",
  1868 => x"e2b00c73",
  1869 => x"8f0680e2",
  1870 => x"ac0ca052",
  1871 => x"7380e380",
  1872 => x"082e0981",
  1873 => x"06993880",
  1874 => x"e2fc08ff",
  1875 => x"05743270",
  1876 => x"09810570",
  1877 => x"72079f2a",
  1878 => x"91713151",
  1879 => x"51535371",
  1880 => x"5183842d",
  1881 => x"8114548e",
  1882 => x"7425c238",
  1883 => x"80e0b008",
  1884 => x"527180e2",
  1885 => x"9c0c0298",
  1886 => x"050d0402",
  1887 => x"f4050dd4",
  1888 => x"5281ff72",
  1889 => x"0c710853",
  1890 => x"81ff720c",
  1891 => x"72882b83",
  1892 => x"fe800672",
  1893 => x"087081ff",
  1894 => x"06515253",
  1895 => x"81ff720c",
  1896 => x"72710788",
  1897 => x"2b720870",
  1898 => x"81ff0651",
  1899 => x"525381ff",
  1900 => x"720c7271",
  1901 => x"07882b72",
  1902 => x"087081ff",
  1903 => x"06720780",
  1904 => x"e29c0c52",
  1905 => x"53028c05",
  1906 => x"0d0402f4",
  1907 => x"050d7476",
  1908 => x"7181ff06",
  1909 => x"d40c5353",
  1910 => x"80e38808",
  1911 => x"85387189",
  1912 => x"2b527198",
  1913 => x"2ad40c71",
  1914 => x"902a7081",
  1915 => x"ff06d40c",
  1916 => x"5171882a",
  1917 => x"7081ff06",
  1918 => x"d40c5171",
  1919 => x"81ff06d4",
  1920 => x"0c72902a",
  1921 => x"7081ff06",
  1922 => x"d40c51d4",
  1923 => x"087081ff",
  1924 => x"06515182",
  1925 => x"b8bf5270",
  1926 => x"81ff2e09",
  1927 => x"81069438",
  1928 => x"81ff0bd4",
  1929 => x"0cd40870",
  1930 => x"81ff06ff",
  1931 => x"14545151",
  1932 => x"71e53870",
  1933 => x"80e29c0c",
  1934 => x"028c050d",
  1935 => x"0402fc05",
  1936 => x"0d81c751",
  1937 => x"81ff0bd4",
  1938 => x"0cff1151",
  1939 => x"708025f4",
  1940 => x"38028405",
  1941 => x"0d0402f4",
  1942 => x"050d81ff",
  1943 => x"0bd40c93",
  1944 => x"53805287",
  1945 => x"fc80c151",
  1946 => x"bbca2d80",
  1947 => x"e29c088b",
  1948 => x"3881ff0b",
  1949 => x"d40c8153",
  1950 => x"bd8404bc",
  1951 => x"bd2dff13",
  1952 => x"5372de38",
  1953 => x"7280e29c",
  1954 => x"0c028c05",
  1955 => x"0d0402ec",
  1956 => x"050d810b",
  1957 => x"80e3880c",
  1958 => x"8454d008",
  1959 => x"708f2a70",
  1960 => x"81065151",
  1961 => x"5372f338",
  1962 => x"72d00cbc",
  1963 => x"bd2d80db",
  1964 => x"dc5186a0",
  1965 => x"2dd00870",
  1966 => x"8f2a7081",
  1967 => x"06515153",
  1968 => x"72f33881",
  1969 => x"0bd00cb1",
  1970 => x"53805284",
  1971 => x"d480c051",
  1972 => x"bbca2d80",
  1973 => x"e29c0881",
  1974 => x"2e933872",
  1975 => x"822ebf38",
  1976 => x"ff135372",
  1977 => x"e438ff14",
  1978 => x"5473ffae",
  1979 => x"38bcbd2d",
  1980 => x"83aa5284",
  1981 => x"9c80c851",
  1982 => x"bbca2d80",
  1983 => x"e29c0881",
  1984 => x"2e098106",
  1985 => x"9338bafb",
  1986 => x"2d80e29c",
  1987 => x"0883ffff",
  1988 => x"06537283",
  1989 => x"aa2ea038",
  1990 => x"bcd62dbe",
  1991 => x"b20480db",
  1992 => x"e85186a0",
  1993 => x"2d805380",
  1994 => x"c0870480",
  1995 => x"dc805186",
  1996 => x"a02d8054",
  1997 => x"bfd80481",
  1998 => x"ff0bd40c",
  1999 => x"b154bcbd",
  2000 => x"2d8fcf53",
  2001 => x"805287fc",
  2002 => x"80f751bb",
  2003 => x"ca2d80e2",
  2004 => x"9c085580",
  2005 => x"e29c0881",
  2006 => x"2e098106",
  2007 => x"9c3881ff",
  2008 => x"0bd40c82",
  2009 => x"0a52849c",
  2010 => x"80e951bb",
  2011 => x"ca2d80e2",
  2012 => x"9c08802e",
  2013 => x"8d38bcbd",
  2014 => x"2dff1353",
  2015 => x"72c638bf",
  2016 => x"cb0481ff",
  2017 => x"0bd40c80",
  2018 => x"e29c0852",
  2019 => x"87fc80fa",
  2020 => x"51bbca2d",
  2021 => x"80e29c08",
  2022 => x"b23881ff",
  2023 => x"0bd40cd4",
  2024 => x"085381ff",
  2025 => x"0bd40c81",
  2026 => x"ff0bd40c",
  2027 => x"81ff0bd4",
  2028 => x"0c81ff0b",
  2029 => x"d40c7286",
  2030 => x"2a708106",
  2031 => x"76565153",
  2032 => x"72963880",
  2033 => x"e29c0854",
  2034 => x"bfd80473",
  2035 => x"822efedb",
  2036 => x"38ff1454",
  2037 => x"73fee738",
  2038 => x"7380e388",
  2039 => x"0c738b38",
  2040 => x"815287fc",
  2041 => x"80d051bb",
  2042 => x"ca2d81ff",
  2043 => x"0bd40cd0",
  2044 => x"08708f2a",
  2045 => x"70810651",
  2046 => x"515372f3",
  2047 => x"3872d00c",
  2048 => x"81ff0bd4",
  2049 => x"0c815372",
  2050 => x"80e29c0c",
  2051 => x"0294050d",
  2052 => x"0402e805",
  2053 => x"0d785580",
  2054 => x"5681ff0b",
  2055 => x"d40cd008",
  2056 => x"708f2a70",
  2057 => x"81065151",
  2058 => x"5372f338",
  2059 => x"82810bd0",
  2060 => x"0c81ff0b",
  2061 => x"d40c7752",
  2062 => x"87fc80d1",
  2063 => x"51bbca2d",
  2064 => x"80dbc6df",
  2065 => x"5480e29c",
  2066 => x"08802e8c",
  2067 => x"3880dca0",
  2068 => x"5186a02d",
  2069 => x"80c1ad04",
  2070 => x"81ff0bd4",
  2071 => x"0cd40870",
  2072 => x"81ff0651",
  2073 => x"537281fe",
  2074 => x"2e098106",
  2075 => x"9f3880ff",
  2076 => x"53bafb2d",
  2077 => x"80e29c08",
  2078 => x"75708405",
  2079 => x"570cff13",
  2080 => x"53728025",
  2081 => x"ec388156",
  2082 => x"80c19204",
  2083 => x"ff145473",
  2084 => x"c73881ff",
  2085 => x"0bd40c81",
  2086 => x"ff0bd40c",
  2087 => x"d008708f",
  2088 => x"2a708106",
  2089 => x"51515372",
  2090 => x"f33872d0",
  2091 => x"0c7580e2",
  2092 => x"9c0c0298",
  2093 => x"050d0402",
  2094 => x"e8050d77",
  2095 => x"797b5855",
  2096 => x"55805372",
  2097 => x"7625a538",
  2098 => x"74708105",
  2099 => x"5680f52d",
  2100 => x"74708105",
  2101 => x"5680f52d",
  2102 => x"52527171",
  2103 => x"2e873881",
  2104 => x"5180c1ee",
  2105 => x"04811353",
  2106 => x"80c1c304",
  2107 => x"80517080",
  2108 => x"e29c0c02",
  2109 => x"98050d04",
  2110 => x"02ec050d",
  2111 => x"7680e9c8",
  2112 => x"55559f53",
  2113 => x"80747084",
  2114 => x"05560cff",
  2115 => x"13537280",
  2116 => x"25f23874",
  2117 => x"802e80c4",
  2118 => x"389a1580",
  2119 => x"e02d5180",
  2120 => x"d2902d80",
  2121 => x"e29c0880",
  2122 => x"e29c0880",
  2123 => x"e9bc0c80",
  2124 => x"e29c0854",
  2125 => x"5480e998",
  2126 => x"08802e9b",
  2127 => x"38941580",
  2128 => x"e02d5180",
  2129 => x"d2902d80",
  2130 => x"e29c0890",
  2131 => x"2b83fff0",
  2132 => x"0a067075",
  2133 => x"07515372",
  2134 => x"80e9bc0c",
  2135 => x"80e9bc08",
  2136 => x"5372802e",
  2137 => x"9e3880e9",
  2138 => x"9008fe14",
  2139 => x"712980e9",
  2140 => x"a4080580",
  2141 => x"e9c00c70",
  2142 => x"842b80e9",
  2143 => x"9c0c5480",
  2144 => x"c3b20480",
  2145 => x"e9a80880",
  2146 => x"e9bc0c80",
  2147 => x"e9ac0880",
  2148 => x"e9c00c80",
  2149 => x"e9980880",
  2150 => x"2e8c3880",
  2151 => x"e9900884",
  2152 => x"2b5380c3",
  2153 => x"ad0480e9",
  2154 => x"b008842b",
  2155 => x"537280e9",
  2156 => x"9c0c0294",
  2157 => x"050d0402",
  2158 => x"d8050d80",
  2159 => x"0b80e998",
  2160 => x"0c8454bd",
  2161 => x"8e2d80e2",
  2162 => x"9c08802e",
  2163 => x"993880e3",
  2164 => x"8c528051",
  2165 => x"80c0912d",
  2166 => x"80e29c08",
  2167 => x"802e8738",
  2168 => x"fe5480c3",
  2169 => x"ee04ff14",
  2170 => x"54738024",
  2171 => x"d638738e",
  2172 => x"3880dcb0",
  2173 => x"5186a02d",
  2174 => x"735580c9",
  2175 => x"d2048056",
  2176 => x"810b80e9",
  2177 => x"c40c8853",
  2178 => x"80dcc452",
  2179 => x"80e3c251",
  2180 => x"80c1b72d",
  2181 => x"80e29c08",
  2182 => x"762e0981",
  2183 => x"06893880",
  2184 => x"e29c0880",
  2185 => x"e9c40c88",
  2186 => x"5380dcd0",
  2187 => x"5280e3de",
  2188 => x"5180c1b7",
  2189 => x"2d80e29c",
  2190 => x"08893880",
  2191 => x"e29c0880",
  2192 => x"e9c40c80",
  2193 => x"e9c40880",
  2194 => x"2e818538",
  2195 => x"80e6d20b",
  2196 => x"80f52d80",
  2197 => x"e6d30b80",
  2198 => x"f52d7198",
  2199 => x"2b71902b",
  2200 => x"0780e6d4",
  2201 => x"0b80f52d",
  2202 => x"70882b72",
  2203 => x"0780e6d5",
  2204 => x"0b80f52d",
  2205 => x"710780e7",
  2206 => x"8a0b80f5",
  2207 => x"2d80e78b",
  2208 => x"0b80f52d",
  2209 => x"71882b07",
  2210 => x"535f5452",
  2211 => x"5a565755",
  2212 => x"7381abaa",
  2213 => x"2e098106",
  2214 => x"90387551",
  2215 => x"80d1df2d",
  2216 => x"80e29c08",
  2217 => x"5680c5b8",
  2218 => x"047382d4",
  2219 => x"d52e8938",
  2220 => x"80dcdc51",
  2221 => x"80c68804",
  2222 => x"80e38c52",
  2223 => x"755180c0",
  2224 => x"912d80e2",
  2225 => x"9c085580",
  2226 => x"e29c0880",
  2227 => x"2e848338",
  2228 => x"885380dc",
  2229 => x"d05280e3",
  2230 => x"de5180c1",
  2231 => x"b72d80e2",
  2232 => x"9c088b38",
  2233 => x"810b80e9",
  2234 => x"980c80c6",
  2235 => x"8f048853",
  2236 => x"80dcc452",
  2237 => x"80e3c251",
  2238 => x"80c1b72d",
  2239 => x"80e29c08",
  2240 => x"802e8c38",
  2241 => x"80dcf051",
  2242 => x"86a02d80",
  2243 => x"c6ee0480",
  2244 => x"e78a0b80",
  2245 => x"f52d5473",
  2246 => x"80d52e09",
  2247 => x"810680ce",
  2248 => x"3880e78b",
  2249 => x"0b80f52d",
  2250 => x"547381aa",
  2251 => x"2e098106",
  2252 => x"bd38800b",
  2253 => x"80e38c0b",
  2254 => x"80f52d56",
  2255 => x"547481e9",
  2256 => x"2e833881",
  2257 => x"547481eb",
  2258 => x"2e8c3880",
  2259 => x"5573752e",
  2260 => x"09810682",
  2261 => x"fd3880e3",
  2262 => x"970b80f5",
  2263 => x"2d55748e",
  2264 => x"3880e398",
  2265 => x"0b80f52d",
  2266 => x"5473822e",
  2267 => x"87388055",
  2268 => x"80c9d204",
  2269 => x"80e3990b",
  2270 => x"80f52d70",
  2271 => x"80e9900c",
  2272 => x"ff0580e9",
  2273 => x"940c80e3",
  2274 => x"9a0b80f5",
  2275 => x"2d80e39b",
  2276 => x"0b80f52d",
  2277 => x"58760577",
  2278 => x"82802905",
  2279 => x"7080e9a0",
  2280 => x"0c80e39c",
  2281 => x"0b80f52d",
  2282 => x"7080e9b4",
  2283 => x"0c80e998",
  2284 => x"08595758",
  2285 => x"76802e81",
  2286 => x"b9388853",
  2287 => x"80dcd052",
  2288 => x"80e3de51",
  2289 => x"80c1b72d",
  2290 => x"80e29c08",
  2291 => x"82843880",
  2292 => x"e9900870",
  2293 => x"842b80e9",
  2294 => x"9c0c7080",
  2295 => x"e9b00c80",
  2296 => x"e3b10b80",
  2297 => x"f52d80e3",
  2298 => x"b00b80f5",
  2299 => x"2d718280",
  2300 => x"290580e3",
  2301 => x"b20b80f5",
  2302 => x"2d708480",
  2303 => x"80291280",
  2304 => x"e3b30b80",
  2305 => x"f52d7081",
  2306 => x"800a2912",
  2307 => x"7080e9b8",
  2308 => x"0c80e9b4",
  2309 => x"08712980",
  2310 => x"e9a00805",
  2311 => x"7080e9a4",
  2312 => x"0c80e3b9",
  2313 => x"0b80f52d",
  2314 => x"80e3b80b",
  2315 => x"80f52d71",
  2316 => x"82802905",
  2317 => x"80e3ba0b",
  2318 => x"80f52d70",
  2319 => x"84808029",
  2320 => x"1280e3bb",
  2321 => x"0b80f52d",
  2322 => x"70982b81",
  2323 => x"f00a0672",
  2324 => x"057080e9",
  2325 => x"a80cfe11",
  2326 => x"7e297705",
  2327 => x"80e9ac0c",
  2328 => x"52595243",
  2329 => x"545e5152",
  2330 => x"59525d57",
  2331 => x"595780c9",
  2332 => x"ca0480e3",
  2333 => x"9e0b80f5",
  2334 => x"2d80e39d",
  2335 => x"0b80f52d",
  2336 => x"71828029",
  2337 => x"057080e9",
  2338 => x"9c0c70a0",
  2339 => x"2983ff05",
  2340 => x"70892a70",
  2341 => x"80e9b00c",
  2342 => x"80e3a30b",
  2343 => x"80f52d80",
  2344 => x"e3a20b80",
  2345 => x"f52d7182",
  2346 => x"80290570",
  2347 => x"80e9b80c",
  2348 => x"7b71291e",
  2349 => x"7080e9ac",
  2350 => x"0c7d80e9",
  2351 => x"a80c7305",
  2352 => x"80e9a40c",
  2353 => x"555e5151",
  2354 => x"55558051",
  2355 => x"80c1f82d",
  2356 => x"81557480",
  2357 => x"e29c0c02",
  2358 => x"a8050d04",
  2359 => x"02ec050d",
  2360 => x"7670872c",
  2361 => x"7180ff06",
  2362 => x"55565480",
  2363 => x"e998088a",
  2364 => x"3873882c",
  2365 => x"7481ff06",
  2366 => x"545580e3",
  2367 => x"8c5280e9",
  2368 => x"a0081551",
  2369 => x"80c0912d",
  2370 => x"80e29c08",
  2371 => x"5480e29c",
  2372 => x"08802ebb",
  2373 => x"3880e998",
  2374 => x"08802e9c",
  2375 => x"38728429",
  2376 => x"80e38c05",
  2377 => x"70085253",
  2378 => x"80d1df2d",
  2379 => x"80e29c08",
  2380 => x"f00a0653",
  2381 => x"80cacd04",
  2382 => x"721080e3",
  2383 => x"8c057080",
  2384 => x"e02d5253",
  2385 => x"80d2902d",
  2386 => x"80e29c08",
  2387 => x"53725473",
  2388 => x"80e29c0c",
  2389 => x"0294050d",
  2390 => x"0402dc05",
  2391 => x"0d7a7c59",
  2392 => x"55805477",
  2393 => x"742e8438",
  2394 => x"73780c74",
  2395 => x"842c80e9",
  2396 => x"c0080575",
  2397 => x"8f065459",
  2398 => x"7281a038",
  2399 => x"80e99808",
  2400 => x"802e818d",
  2401 => x"3880e9bc",
  2402 => x"085680e9",
  2403 => x"9c087526",
  2404 => x"80f73880",
  2405 => x"e9c85773",
  2406 => x"9f268f38",
  2407 => x"76085372",
  2408 => x"802e8738",
  2409 => x"725680cb",
  2410 => x"d5047551",
  2411 => x"80c9dc2d",
  2412 => x"80e29c08",
  2413 => x"80e29c08",
  2414 => x"80ffffff",
  2415 => x"f8065456",
  2416 => x"7280ffff",
  2417 => x"fff82e83",
  2418 => x"8a38739f",
  2419 => x"26873880",
  2420 => x"e29c0877",
  2421 => x"0c80e99c",
  2422 => x"08757131",
  2423 => x"8116841a",
  2424 => x"5a565653",
  2425 => x"747327ff",
  2426 => x"ae387380",
  2427 => x"2e9b38fe",
  2428 => x"1680e990",
  2429 => x"082980e9",
  2430 => x"a4080575",
  2431 => x"842c0576",
  2432 => x"80e0b40c",
  2433 => x"5980cc91",
  2434 => x"0480e9bc",
  2435 => x"0880e0b4",
  2436 => x"0c80e38c",
  2437 => x"52785180",
  2438 => x"c0912d74",
  2439 => x"852b83e0",
  2440 => x"0680e38c",
  2441 => x"05548074",
  2442 => x"80f52d54",
  2443 => x"5672762e",
  2444 => x"09810683",
  2445 => x"38815677",
  2446 => x"802e8f38",
  2447 => x"81707706",
  2448 => x"54557280",
  2449 => x"2e843874",
  2450 => x"780c8074",
  2451 => x"80f52d56",
  2452 => x"5374732e",
  2453 => x"83388153",
  2454 => x"7481e52e",
  2455 => x"81f53881",
  2456 => x"70740654",
  2457 => x"5872802e",
  2458 => x"81e9388b",
  2459 => x"1480f52d",
  2460 => x"70832a79",
  2461 => x"06585676",
  2462 => x"9c3880e0",
  2463 => x"b8085372",
  2464 => x"89387280",
  2465 => x"e78c0b81",
  2466 => x"b72d7680",
  2467 => x"e0b80c73",
  2468 => x"5380ced5",
  2469 => x"04758f2e",
  2470 => x"09810681",
  2471 => x"b638749f",
  2472 => x"068d2980",
  2473 => x"e6ff1151",
  2474 => x"53811480",
  2475 => x"f52d7370",
  2476 => x"81055581",
  2477 => x"b72d8314",
  2478 => x"80f52d73",
  2479 => x"70810555",
  2480 => x"81b72d85",
  2481 => x"1480f52d",
  2482 => x"73708105",
  2483 => x"5581b72d",
  2484 => x"871480f5",
  2485 => x"2d737081",
  2486 => x"055581b7",
  2487 => x"2d891480",
  2488 => x"f52d7370",
  2489 => x"81055581",
  2490 => x"b72d8e14",
  2491 => x"80f52d73",
  2492 => x"70810555",
  2493 => x"81b72d90",
  2494 => x"1480f52d",
  2495 => x"73708105",
  2496 => x"5581b72d",
  2497 => x"921480f5",
  2498 => x"2d737081",
  2499 => x"055581b7",
  2500 => x"2d941480",
  2501 => x"f52d7370",
  2502 => x"81055581",
  2503 => x"b72d9614",
  2504 => x"80f52d73",
  2505 => x"70810555",
  2506 => x"81b72d98",
  2507 => x"1480f52d",
  2508 => x"73708105",
  2509 => x"5581b72d",
  2510 => x"9c1480f5",
  2511 => x"2d737081",
  2512 => x"055581b7",
  2513 => x"2d9e1480",
  2514 => x"f52d7381",
  2515 => x"b72d7780",
  2516 => x"e0b80c80",
  2517 => x"537280e2",
  2518 => x"9c0c02a4",
  2519 => x"050d0402",
  2520 => x"cc050d7e",
  2521 => x"605e5a80",
  2522 => x"0b80e9bc",
  2523 => x"0880e9c0",
  2524 => x"08595c56",
  2525 => x"805880e9",
  2526 => x"9c08782e",
  2527 => x"81be3877",
  2528 => x"8f06a017",
  2529 => x"57547392",
  2530 => x"3880e38c",
  2531 => x"52765181",
  2532 => x"175780c0",
  2533 => x"912d80e3",
  2534 => x"8c568076",
  2535 => x"80f52d56",
  2536 => x"5474742e",
  2537 => x"83388154",
  2538 => x"7481e52e",
  2539 => x"81823881",
  2540 => x"70750655",
  2541 => x"5c73802e",
  2542 => x"80f6388b",
  2543 => x"1680f52d",
  2544 => x"98065978",
  2545 => x"80ea388b",
  2546 => x"537c5275",
  2547 => x"5180c1b7",
  2548 => x"2d80e29c",
  2549 => x"0880d938",
  2550 => x"9c160851",
  2551 => x"80d1df2d",
  2552 => x"80e29c08",
  2553 => x"841b0c9a",
  2554 => x"1680e02d",
  2555 => x"5180d290",
  2556 => x"2d80e29c",
  2557 => x"0880e29c",
  2558 => x"08881c0c",
  2559 => x"80e29c08",
  2560 => x"555580e9",
  2561 => x"9808802e",
  2562 => x"9a389416",
  2563 => x"80e02d51",
  2564 => x"80d2902d",
  2565 => x"80e29c08",
  2566 => x"902b83ff",
  2567 => x"f00a0670",
  2568 => x"16515473",
  2569 => x"881b0c78",
  2570 => x"7a0c7b54",
  2571 => x"80d0fa04",
  2572 => x"81185880",
  2573 => x"e99c0878",
  2574 => x"26fec438",
  2575 => x"80e99808",
  2576 => x"802eb538",
  2577 => x"7a5180c9",
  2578 => x"dc2d80e2",
  2579 => x"9c0880e2",
  2580 => x"9c0880ff",
  2581 => x"fffff806",
  2582 => x"555b7380",
  2583 => x"fffffff8",
  2584 => x"2e963880",
  2585 => x"e29c08fe",
  2586 => x"0580e990",
  2587 => x"082980e9",
  2588 => x"a4080557",
  2589 => x"80cef404",
  2590 => x"80547380",
  2591 => x"e29c0c02",
  2592 => x"b4050d04",
  2593 => x"02f4050d",
  2594 => x"74700881",
  2595 => x"05710c70",
  2596 => x"0880e994",
  2597 => x"08065353",
  2598 => x"71903888",
  2599 => x"13085180",
  2600 => x"c9dc2d80",
  2601 => x"e29c0888",
  2602 => x"140c810b",
  2603 => x"80e29c0c",
  2604 => x"028c050d",
  2605 => x"0402f005",
  2606 => x"0d758811",
  2607 => x"08fe0580",
  2608 => x"e9900829",
  2609 => x"80e9a408",
  2610 => x"11720880",
  2611 => x"e9940806",
  2612 => x"05795553",
  2613 => x"545480c0",
  2614 => x"912d0290",
  2615 => x"050d0402",
  2616 => x"f4050d74",
  2617 => x"70882a83",
  2618 => x"fe800670",
  2619 => x"72982a07",
  2620 => x"72882b87",
  2621 => x"fc808006",
  2622 => x"73982b81",
  2623 => x"f00a0671",
  2624 => x"73070780",
  2625 => x"e29c0c56",
  2626 => x"51535102",
  2627 => x"8c050d04",
  2628 => x"02f8050d",
  2629 => x"028e0580",
  2630 => x"f52d7488",
  2631 => x"2b077083",
  2632 => x"ffff0680",
  2633 => x"e29c0c51",
  2634 => x"0288050d",
  2635 => x"0402f405",
  2636 => x"0d747678",
  2637 => x"53545280",
  2638 => x"71259738",
  2639 => x"72708105",
  2640 => x"5480f52d",
  2641 => x"72708105",
  2642 => x"5481b72d",
  2643 => x"ff115170",
  2644 => x"eb388072",
  2645 => x"81b72d02",
  2646 => x"8c050d04",
  2647 => x"02e0050d",
  2648 => x"79578070",
  2649 => x"59705755",
  2650 => x"80d39304",
  2651 => x"02a005fc",
  2652 => x"05527551",
  2653 => x"80cad92d",
  2654 => x"80e29c08",
  2655 => x"80e29c08",
  2656 => x"09810570",
  2657 => x"80e29c08",
  2658 => x"079f2a77",
  2659 => x"05811959",
  2660 => x"57545476",
  2661 => x"75255377",
  2662 => x"843872d0",
  2663 => x"387380e2",
  2664 => x"9c0c02a0",
  2665 => x"050d0402",
  2666 => x"f0050d80",
  2667 => x"e2980816",
  2668 => x"5180d2dc",
  2669 => x"2d80e29c",
  2670 => x"08802ea0",
  2671 => x"388b5380",
  2672 => x"e29c0852",
  2673 => x"80e78c51",
  2674 => x"80d2ad2d",
  2675 => x"80eac808",
  2676 => x"5473802e",
  2677 => x"873880e7",
  2678 => x"8c51732d",
  2679 => x"0290050d",
  2680 => x"0402f405",
  2681 => x"0d747670",
  2682 => x"8c2c708f",
  2683 => x"0680dda0",
  2684 => x"08055153",
  2685 => x"53537080",
  2686 => x"f52d7381",
  2687 => x"b72d7188",
  2688 => x"2c708f06",
  2689 => x"80dda008",
  2690 => x"05515170",
  2691 => x"80f52d81",
  2692 => x"1481b72d",
  2693 => x"71842c70",
  2694 => x"8f0680dd",
  2695 => x"a0080551",
  2696 => x"517080f5",
  2697 => x"2d821481",
  2698 => x"b72d718f",
  2699 => x"0680dda0",
  2700 => x"08055271",
  2701 => x"80f52d83",
  2702 => x"1481b72d",
  2703 => x"028c050d",
  2704 => x"0402d805",
  2705 => x"0d805a80",
  2706 => x"70565980",
  2707 => x"d4f10402",
  2708 => x"a805fc05",
  2709 => x"52785180",
  2710 => x"cad92d80",
  2711 => x"e29c0809",
  2712 => x"81057080",
  2713 => x"e29c0807",
  2714 => x"9f2a7605",
  2715 => x"811b5b56",
  2716 => x"5480e298",
  2717 => x"08752454",
  2718 => x"79843873",
  2719 => x"d2388070",
  2720 => x"5b5502a8",
  2721 => x"05fc0552",
  2722 => x"785180ca",
  2723 => x"d92d80e2",
  2724 => x"9c08802e",
  2725 => x"81b43880",
  2726 => x"e29c088b",
  2727 => x"0580f52d",
  2728 => x"70842a70",
  2729 => x"81067710",
  2730 => x"78842b80",
  2731 => x"e78c0b80",
  2732 => x"f52d5c5c",
  2733 => x"53515556",
  2734 => x"73802e80",
  2735 => x"ce387416",
  2736 => x"822b80d8",
  2737 => x"e00b80e0",
  2738 => x"c4120c54",
  2739 => x"77753110",
  2740 => x"80eacc11",
  2741 => x"55569074",
  2742 => x"70810556",
  2743 => x"81b72da0",
  2744 => x"7481b72d",
  2745 => x"7681ff06",
  2746 => x"81165854",
  2747 => x"73802e8b",
  2748 => x"389c5380",
  2749 => x"e78c5280",
  2750 => x"d682048b",
  2751 => x"5380e29c",
  2752 => x"085280ea",
  2753 => x"ce165180",
  2754 => x"d6c00474",
  2755 => x"16822b80",
  2756 => x"d3a70b80",
  2757 => x"e0c4120c",
  2758 => x"547681ff",
  2759 => x"06811658",
  2760 => x"5473802e",
  2761 => x"8b389c53",
  2762 => x"80e78c52",
  2763 => x"80d6b704",
  2764 => x"8b5380e2",
  2765 => x"9c085277",
  2766 => x"75311080",
  2767 => x"eacc0551",
  2768 => x"765580d2",
  2769 => x"ad2d80d6",
  2770 => x"df047490",
  2771 => x"29753170",
  2772 => x"1080eacc",
  2773 => x"05515480",
  2774 => x"e29c0874",
  2775 => x"81b72d81",
  2776 => x"1959748b",
  2777 => x"24a63879",
  2778 => x"802efe96",
  2779 => x"38749029",
  2780 => x"75317010",
  2781 => x"80eacc05",
  2782 => x"8c773157",
  2783 => x"51548074",
  2784 => x"81b72d9e",
  2785 => x"14ff1656",
  2786 => x"5474f338",
  2787 => x"80dcfc52",
  2788 => x"80e1f051",
  2789 => x"a2ce2d80",
  2790 => x"e2980852",
  2791 => x"80e1f551",
  2792 => x"80d3e12d",
  2793 => x"80e99c08",
  2794 => x"5280e1fa",
  2795 => x"5180d3e1",
  2796 => x"2d785280",
  2797 => x"e1ff5180",
  2798 => x"d3e12d80",
  2799 => x"e0b40b80",
  2800 => x"e02d5280",
  2801 => x"e2845180",
  2802 => x"d3e12d80",
  2803 => x"e0b60b80",
  2804 => x"e02d5280",
  2805 => x"e2885180",
  2806 => x"d3e12d78",
  2807 => x"80e29c0c",
  2808 => x"02a8050d",
  2809 => x"0402fc05",
  2810 => x"0d725170",
  2811 => x"fd2eb238",
  2812 => x"70fd248b",
  2813 => x"3870fc2e",
  2814 => x"80d03880",
  2815 => x"d8d40470",
  2816 => x"fe2eb938",
  2817 => x"70ff2e09",
  2818 => x"810680c8",
  2819 => x"3880e298",
  2820 => x"08517080",
  2821 => x"2ebe38ff",
  2822 => x"1180e298",
  2823 => x"0c80d8d4",
  2824 => x"0480e298",
  2825 => x"08f40570",
  2826 => x"80e2980c",
  2827 => x"51708025",
  2828 => x"a338800b",
  2829 => x"80e2980c",
  2830 => x"80d8d404",
  2831 => x"80e29808",
  2832 => x"810580e2",
  2833 => x"980c80d8",
  2834 => x"d40480e2",
  2835 => x"98088c05",
  2836 => x"80e2980c",
  2837 => x"80d4c12d",
  2838 => x"affd2d02",
  2839 => x"84050d04",
  2840 => x"02fc050d",
  2841 => x"80e29808",
  2842 => x"135180d2",
  2843 => x"dc2d80e2",
  2844 => x"9c08802e",
  2845 => x"8a3880e2",
  2846 => x"9c085180",
  2847 => x"c1f82d80",
  2848 => x"0b80e298",
  2849 => x"0c80d4c1",
  2850 => x"2daffd2d",
  2851 => x"0284050d",
  2852 => x"0402fc05",
  2853 => x"0d800b80",
  2854 => x"e2980c80",
  2855 => x"d4c12dae",
  2856 => x"f92d80e2",
  2857 => x"9c0880e1",
  2858 => x"e00c80e0",
  2859 => x"bc51b1a3",
  2860 => x"2d028405",
  2861 => x"0d047180",
  2862 => x"eac80c04",
  2863 => x"00ffffff",
  2864 => x"ff00ffff",
  2865 => x"ffff00ff",
  2866 => x"ffffff00",
  2867 => x"30313233",
  2868 => x"34353637",
  2869 => x"38394142",
  2870 => x"43444546",
  2871 => x"00000000",
  2872 => x"52657365",
  2873 => x"74000000",
  2874 => x"5363616e",
  2875 => x"6c696e65",
  2876 => x"73000000",
  2877 => x"50414c20",
  2878 => x"2f204e54",
  2879 => x"53430000",
  2880 => x"436f6c6f",
  2881 => x"72000000",
  2882 => x"44696666",
  2883 => x"6963756c",
  2884 => x"74792041",
  2885 => x"00000000",
  2886 => x"44696666",
  2887 => x"6963756c",
  2888 => x"74792042",
  2889 => x"00000000",
  2890 => x"2a537570",
  2891 => x"65726368",
  2892 => x"69702069",
  2893 => x"6e206361",
  2894 => x"72747269",
  2895 => x"64676500",
  2896 => x"2a42616e",
  2897 => x"6b204530",
  2898 => x"00000000",
  2899 => x"2a42616e",
  2900 => x"6b204537",
  2901 => x"00000000",
  2902 => x"53656c65",
  2903 => x"63740000",
  2904 => x"53746172",
  2905 => x"74000000",
  2906 => x"4c6f6164",
  2907 => x"20524f4d",
  2908 => x"20100000",
  2909 => x"45786974",
  2910 => x"00000000",
  2911 => x"43617274",
  2912 => x"72696467",
  2913 => x"65000000",
  2914 => x"524f4d20",
  2915 => x"6c6f6164",
  2916 => x"696e6720",
  2917 => x"6661696c",
  2918 => x"65640000",
  2919 => x"4f4b0000",
  2920 => x"496e6974",
  2921 => x"69616c69",
  2922 => x"7a696e67",
  2923 => x"20534420",
  2924 => x"63617264",
  2925 => x"0a000000",
  2926 => x"446f6e65",
  2927 => x"20696e69",
  2928 => x"7469616c",
  2929 => x"697a6174",
  2930 => x"696f6e0a",
  2931 => x"00000000",
  2932 => x"16200000",
  2933 => x"14200000",
  2934 => x"15200000",
  2935 => x"53442069",
  2936 => x"6e69742e",
  2937 => x"2e2e0a00",
  2938 => x"53442063",
  2939 => x"61726420",
  2940 => x"72657365",
  2941 => x"74206661",
  2942 => x"696c6564",
  2943 => x"210a0000",
  2944 => x"53444843",
  2945 => x"20657272",
  2946 => x"6f72210a",
  2947 => x"00000000",
  2948 => x"57726974",
  2949 => x"65206661",
  2950 => x"696c6564",
  2951 => x"0a000000",
  2952 => x"52656164",
  2953 => x"20666169",
  2954 => x"6c65640a",
  2955 => x"00000000",
  2956 => x"43617264",
  2957 => x"20696e69",
  2958 => x"74206661",
  2959 => x"696c6564",
  2960 => x"0a000000",
  2961 => x"46415431",
  2962 => x"36202020",
  2963 => x"00000000",
  2964 => x"46415433",
  2965 => x"32202020",
  2966 => x"00000000",
  2967 => x"4e6f2070",
  2968 => x"61727469",
  2969 => x"74696f6e",
  2970 => x"20736967",
  2971 => x"0a000000",
  2972 => x"42616420",
  2973 => x"70617274",
  2974 => x"0a000000",
  2975 => x"4261636b",
  2976 => x"20787878",
  2977 => x"78207979",
  2978 => x"7979207a",
  2979 => x"7a7a7a20",
  2980 => x"6b6b6b6b",
  2981 => x"6b6b6b6b",
  2982 => x"00000000",
  2983 => x"00000002",
  2984 => x"00002ccc",
  2985 => x"00000002",
  2986 => x"00002ce0",
  2987 => x"0000035a",
  2988 => x"00000001",
  2989 => x"00002ce8",
  2990 => x"00000000",
  2991 => x"00000001",
  2992 => x"00002cf4",
  2993 => x"00000001",
  2994 => x"00000001",
  2995 => x"00002d00",
  2996 => x"00000002",
  2997 => x"00000001",
  2998 => x"00002d08",
  2999 => x"00000003",
  3000 => x"00000001",
  3001 => x"00002d18",
  3002 => x"00000004",
  3003 => x"00000001",
  3004 => x"00002d28",
  3005 => x"00000005",
  3006 => x"00000001",
  3007 => x"00002d40",
  3008 => x"00000008",
  3009 => x"00000001",
  3010 => x"00002d4c",
  3011 => x"00000009",
  3012 => x"00000002",
  3013 => x"00002d58",
  3014 => x"0000036e",
  3015 => x"00000002",
  3016 => x"00002d60",
  3017 => x"00000a3f",
  3018 => x"00000002",
  3019 => x"00002d68",
  3020 => x"00002c91",
  3021 => x"00000002",
  3022 => x"00002d74",
  3023 => x"00001796",
  3024 => x"00000002",
  3025 => x"00002d7c",
  3026 => x"00001124",
  3027 => x"00000000",
  3028 => x"00000000",
  3029 => x"00000000",
  3030 => x"00000004",
  3031 => x"00002d88",
  3032 => x"00002f58",
  3033 => x"00000004",
  3034 => x"00002d9c",
  3035 => x"00002ea4",
  3036 => x"00000000",
  3037 => x"00000000",
  3038 => x"00000000",
  3039 => x"00000000",
  3040 => x"00000000",
  3041 => x"00000000",
  3042 => x"00000000",
  3043 => x"00000000",
  3044 => x"00000000",
  3045 => x"00000000",
  3046 => x"00000000",
  3047 => x"00000000",
  3048 => x"00000000",
  3049 => x"00000000",
  3050 => x"00000000",
  3051 => x"00000000",
  3052 => x"00000000",
  3053 => x"00000000",
  3054 => x"00000000",
  3055 => x"761c1c1c",
  3056 => x"1c1c051c",
  3057 => x"1c1c1c1c",
  3058 => x"f2f5fafd",
  3059 => x"5a000000",
  3060 => x"00000000",
  3061 => x"00000000",
  3062 => x"00000000",
  3063 => x"00000000",
  3064 => x"00000000",
  3065 => x"00000000",
  3066 => x"00000000",
  3067 => x"00000000",
  3068 => x"00000000",
  3069 => x"00000000",
  3070 => x"00000000",
  3071 => x"00000000",
  3072 => x"00000000",
  3073 => x"00000000",
  3074 => x"00000000",
  3075 => x"00000000",
  3076 => x"00000000",
  3077 => x"00000000",
  3078 => x"0001ffff",
  3079 => x"0001ffff",
  3080 => x"0001ffff",
  3081 => x"00000000",
  3082 => x"00000000",
  3083 => x"00000004",
  3084 => x"00000000",
  3085 => x"00000000",
  3086 => x"00000000",
  3087 => x"00000002",
  3088 => x"0000354c",
  3089 => x"000029a7",
  3090 => x"00000002",
  3091 => x"0000356a",
  3092 => x"000029a7",
  3093 => x"00000002",
  3094 => x"00003588",
  3095 => x"000029a7",
  3096 => x"00000002",
  3097 => x"000035a6",
  3098 => x"000029a7",
  3099 => x"00000002",
  3100 => x"000035c4",
  3101 => x"000029a7",
  3102 => x"00000002",
  3103 => x"000035e2",
  3104 => x"000029a7",
  3105 => x"00000002",
  3106 => x"00003600",
  3107 => x"000029a7",
  3108 => x"00000002",
  3109 => x"0000361e",
  3110 => x"000029a7",
  3111 => x"00000002",
  3112 => x"0000363c",
  3113 => x"000029a7",
  3114 => x"00000002",
  3115 => x"0000365a",
  3116 => x"000029a7",
  3117 => x"00000002",
  3118 => x"00003678",
  3119 => x"000029a7",
  3120 => x"00000002",
  3121 => x"00003696",
  3122 => x"000029a7",
  3123 => x"00000002",
  3124 => x"000036b4",
  3125 => x"000029a7",
  3126 => x"00000004",
  3127 => x"000030f0",
  3128 => x"00000000",
  3129 => x"00000000",
  3130 => x"00000000",
  3131 => x"00002be5",
  3132 => x"4261636b",
  3133 => x"00000000",
  3134 => x"00000000",
  3135 => x"00000000",
  3136 => x"00000000",
  3137 => x"00000000",
  3138 => x"00000000",
  3139 => x"00000000",
  3140 => x"00000000",
  3141 => x"00000000",
  3142 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

