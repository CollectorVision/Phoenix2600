-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80e1",
     9 => x"80080b0b",
    10 => x"80e18408",
    11 => x"0b0b80e1",
    12 => x"88080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"e1880c0b",
    16 => x"0b80e184",
    17 => x"0c0b0b80",
    18 => x"e1800c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d8dc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80e18070",
    57 => x"80ed8427",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a9b5",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80e1",
    65 => x"900c9f0b",
    66 => x"80e1940c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"e19408ff",
    70 => x"0580e194",
    71 => x"0c80e194",
    72 => x"088025e8",
    73 => x"3880e190",
    74 => x"08ff0580",
    75 => x"e1900c80",
    76 => x"e1900880",
    77 => x"25d03880",
    78 => x"0b80e194",
    79 => x"0c800b80",
    80 => x"e1900c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80e19008",
   100 => x"25913882",
   101 => x"c82d80e1",
   102 => x"9008ff05",
   103 => x"80e1900c",
   104 => x"838a0480",
   105 => x"e1900880",
   106 => x"e1940853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80e19008",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"e1940881",
   116 => x"0580e194",
   117 => x"0c80e194",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80e194",
   121 => x"0c80e190",
   122 => x"08810580",
   123 => x"e1900c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480e1",
   128 => x"94088105",
   129 => x"80e1940c",
   130 => x"80e19408",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80e194",
   134 => x"0c80e190",
   135 => x"08810580",
   136 => x"e1900c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"e1980cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"e1980c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280e1",
   177 => x"98088407",
   178 => x"80e1980c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80dc",
   183 => x"980c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80e198",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80e1",
   208 => x"800c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02f8050d",
  1093 => x"028f0580",
  1094 => x"f52d80dc",
  1095 => x"a0085252",
  1096 => x"7080e2f1",
  1097 => x"279a3871",
  1098 => x"7181b72d",
  1099 => x"80dca008",
  1100 => x"810580dc",
  1101 => x"a00c80dc",
  1102 => x"a0085180",
  1103 => x"7181b72d",
  1104 => x"0288050d",
  1105 => x"0402f405",
  1106 => x"0d747084",
  1107 => x"2a708f06",
  1108 => x"80dc9c08",
  1109 => x"057080f5",
  1110 => x"2d545153",
  1111 => x"53a2902d",
  1112 => x"728f0680",
  1113 => x"dc9c0805",
  1114 => x"7080f52d",
  1115 => x"5253a290",
  1116 => x"2d028c05",
  1117 => x"0d0402f4",
  1118 => x"050d7476",
  1119 => x"54527270",
  1120 => x"81055480",
  1121 => x"f52d5170",
  1122 => x"72708105",
  1123 => x"5481b72d",
  1124 => x"70ec3870",
  1125 => x"7281b72d",
  1126 => x"028c050d",
  1127 => x"0402cc05",
  1128 => x"0d7e5b80",
  1129 => x"0b80dfbc",
  1130 => x"08818006",
  1131 => x"715c5e5c",
  1132 => x"810bec0c",
  1133 => x"840bec0c",
  1134 => x"7a5280e1",
  1135 => x"9c5180cf",
  1136 => x"a62d80e1",
  1137 => x"80087c2e",
  1138 => x"80ff3880",
  1139 => x"e1a0087c",
  1140 => x"ff125759",
  1141 => x"57747c2e",
  1142 => x"8b388118",
  1143 => x"75812a56",
  1144 => x"5874f738",
  1145 => x"f7185881",
  1146 => x"5c807725",
  1147 => x"80db3877",
  1148 => x"52745184",
  1149 => x"a82d80e3",
  1150 => x"bc5280e1",
  1151 => x"9c5180d1",
  1152 => x"fc2d80e1",
  1153 => x"8008802e",
  1154 => x"a63880e3",
  1155 => x"bc597ca7",
  1156 => x"3883ff56",
  1157 => x"78708105",
  1158 => x"5a80f52d",
  1159 => x"7a811c5c",
  1160 => x"e40ce80c",
  1161 => x"ff165675",
  1162 => x"8025e938",
  1163 => x"a4b70480",
  1164 => x"e180085c",
  1165 => x"84805780",
  1166 => x"e19c5180",
  1167 => x"d1cb2dfc",
  1168 => x"80178116",
  1169 => x"5657a3e9",
  1170 => x"0480e1a0",
  1171 => x"08f80c88",
  1172 => x"1b7b5380",
  1173 => x"e1a85255",
  1174 => x"a2f62d80",
  1175 => x"7580f52d",
  1176 => x"7081ff06",
  1177 => x"55585472",
  1178 => x"742eb638",
  1179 => x"811580f5",
  1180 => x"2d537274",
  1181 => x"2eab3873",
  1182 => x"821680f5",
  1183 => x"2d545672",
  1184 => x"80d32e09",
  1185 => x"81068338",
  1186 => x"81567280",
  1187 => x"f3327009",
  1188 => x"81057080",
  1189 => x"25780751",
  1190 => x"51537280",
  1191 => x"2e8338a0",
  1192 => x"54807781",
  1193 => x"ff065456",
  1194 => x"7280c52e",
  1195 => x"09810683",
  1196 => x"38815672",
  1197 => x"80e53270",
  1198 => x"09810570",
  1199 => x"80257807",
  1200 => x"51515372",
  1201 => x"802ea438",
  1202 => x"811580f5",
  1203 => x"2d5372b0",
  1204 => x"2e098106",
  1205 => x"89387382",
  1206 => x"800754a5",
  1207 => x"eb0472b7",
  1208 => x"2e098106",
  1209 => x"86387384",
  1210 => x"80075473",
  1211 => x"802e8e38",
  1212 => x"80dfbc08",
  1213 => x"f9df0674",
  1214 => x"0780dfbc",
  1215 => x"0c810be0",
  1216 => x"0c805186",
  1217 => x"da2d86c7",
  1218 => x"2d7b802e",
  1219 => x"883880dc",
  1220 => x"a451a699",
  1221 => x"0480dde4",
  1222 => x"51b3c32d",
  1223 => x"7b80e180",
  1224 => x"0c02b405",
  1225 => x"0d0402ec",
  1226 => x"050d80e2",
  1227 => x"b00b80dc",
  1228 => x"a00c80e2",
  1229 => x"b0558075",
  1230 => x"81b72d80",
  1231 => x"de880851",
  1232 => x"a2c52dba",
  1233 => x"51a2902d",
  1234 => x"ffb408ff",
  1235 => x"b8087098",
  1236 => x"2a535154",
  1237 => x"a2c52d73",
  1238 => x"902a7081",
  1239 => x"ff065253",
  1240 => x"a2c52d73",
  1241 => x"882a7081",
  1242 => x"ff065253",
  1243 => x"a2c52d73",
  1244 => x"81ff0651",
  1245 => x"a2c52d74",
  1246 => x"5280e1a8",
  1247 => x"51a2f62d",
  1248 => x"7480dca0",
  1249 => x"0c807581",
  1250 => x"b72d80de",
  1251 => x"e0707070",
  1252 => x"84055208",
  1253 => x"535454a2",
  1254 => x"c52d7208",
  1255 => x"51a2c52d",
  1256 => x"88140851",
  1257 => x"a2c52d80",
  1258 => x"dca00853",
  1259 => x"a07381b7",
  1260 => x"2d80dca0",
  1261 => x"08810580",
  1262 => x"dca00c8c",
  1263 => x"140851a2",
  1264 => x"c52d9014",
  1265 => x"0851a2c5",
  1266 => x"2d941408",
  1267 => x"51a2c52d",
  1268 => x"80dca008",
  1269 => x"53a07381",
  1270 => x"b72d80dc",
  1271 => x"a0088105",
  1272 => x"80dca00c",
  1273 => x"98140851",
  1274 => x"a2c52d74",
  1275 => x"5280e1ec",
  1276 => x"51a2f62d",
  1277 => x"80dca451",
  1278 => x"b3c32d80",
  1279 => x"de880884",
  1280 => x"0580de88",
  1281 => x"0c029405",
  1282 => x"0d04800b",
  1283 => x"80de880c",
  1284 => x"0402f405",
  1285 => x"0d80dcb8",
  1286 => x"0b80f52d",
  1287 => x"80dfbc08",
  1288 => x"70810653",
  1289 => x"54527080",
  1290 => x"2e853871",
  1291 => x"84075272",
  1292 => x"812a7081",
  1293 => x"06515170",
  1294 => x"802e8538",
  1295 => x"71820752",
  1296 => x"72822a70",
  1297 => x"81065151",
  1298 => x"70802e85",
  1299 => x"38718107",
  1300 => x"5272832a",
  1301 => x"70810651",
  1302 => x"5170802e",
  1303 => x"85387188",
  1304 => x"07527284",
  1305 => x"2a708106",
  1306 => x"51517080",
  1307 => x"2e853871",
  1308 => x"90075272",
  1309 => x"852a7081",
  1310 => x"06515170",
  1311 => x"802e8538",
  1312 => x"71a00752",
  1313 => x"72882a70",
  1314 => x"81065151",
  1315 => x"70802e86",
  1316 => x"387180c0",
  1317 => x"07527289",
  1318 => x"2a708106",
  1319 => x"51517080",
  1320 => x"2e863871",
  1321 => x"81800752",
  1322 => x"71fc0c71",
  1323 => x"80e1800c",
  1324 => x"028c050d",
  1325 => x"0402f005",
  1326 => x"0d840bec",
  1327 => x"0cb1802d",
  1328 => x"aada2d81",
  1329 => x"f92d8353",
  1330 => x"b0e32d81",
  1331 => x"51858d2d",
  1332 => x"ff135372",
  1333 => x"8025f138",
  1334 => x"840bec0c",
  1335 => x"80dab451",
  1336 => x"86a02d80",
  1337 => x"c5c72d80",
  1338 => x"e1800880",
  1339 => x"2e80d438",
  1340 => x"a39d5180",
  1341 => x"d8d32d80",
  1342 => x"dacc5280",
  1343 => x"e1a851a2",
  1344 => x"f62d80da",
  1345 => x"dc5280e1",
  1346 => x"ec51a2f6",
  1347 => x"2d80dca4",
  1348 => x"51b3c32d",
  1349 => x"b1a22dac",
  1350 => x"852d80e1",
  1351 => x"80088106",
  1352 => x"5372802e",
  1353 => x"86388051",
  1354 => x"94bf2db3",
  1355 => x"d62d80e1",
  1356 => x"800853a8",
  1357 => x"912d8654",
  1358 => x"72833884",
  1359 => x"5473ec0c",
  1360 => x"aa970480",
  1361 => x"0b80e180",
  1362 => x"0c029005",
  1363 => x"0d047198",
  1364 => x"0c04ffb0",
  1365 => x"0880e180",
  1366 => x"0c04810b",
  1367 => x"ffb00c04",
  1368 => x"800bffb0",
  1369 => x"0c0402d8",
  1370 => x"050dffb4",
  1371 => x"0887ffff",
  1372 => x"065a8154",
  1373 => x"807080df",
  1374 => x"a80880df",
  1375 => x"ac0880df",
  1376 => x"845b5957",
  1377 => x"5a587974",
  1378 => x"06757506",
  1379 => x"52527171",
  1380 => x"2e8d3880",
  1381 => x"77818a2d",
  1382 => x"73097506",
  1383 => x"72075576",
  1384 => x"80e02d70",
  1385 => x"83ffff06",
  1386 => x"53517180",
  1387 => x"e42e0981",
  1388 => x"06a23874",
  1389 => x"74067077",
  1390 => x"76063270",
  1391 => x"09810570",
  1392 => x"72079f2a",
  1393 => x"7b057709",
  1394 => x"7a067407",
  1395 => x"5a5b5353",
  1396 => x"53abe204",
  1397 => x"7180e426",
  1398 => x"89388111",
  1399 => x"51707781",
  1400 => x"8a2d7310",
  1401 => x"811a8219",
  1402 => x"595a5490",
  1403 => x"7925ff96",
  1404 => x"387580df",
  1405 => x"ac0c7480",
  1406 => x"dfa80c77",
  1407 => x"80e1800c",
  1408 => x"02a8050d",
  1409 => x"0402d005",
  1410 => x"0d805cad",
  1411 => x"950480e1",
  1412 => x"800881f0",
  1413 => x"2e098106",
  1414 => x"8a38810b",
  1415 => x"80dfb40c",
  1416 => x"ad950480",
  1417 => x"e1800881",
  1418 => x"e02e0981",
  1419 => x"068a3881",
  1420 => x"0b80dfb8",
  1421 => x"0cad9504",
  1422 => x"80e18008",
  1423 => x"5280dfb8",
  1424 => x"08802e89",
  1425 => x"3880e180",
  1426 => x"08818005",
  1427 => x"5271842c",
  1428 => x"728f0653",
  1429 => x"5380dfb4",
  1430 => x"08802e9a",
  1431 => x"38728429",
  1432 => x"80de8c05",
  1433 => x"72138171",
  1434 => x"2b700973",
  1435 => x"0806730c",
  1436 => x"515353ad",
  1437 => x"89047284",
  1438 => x"2980de8c",
  1439 => x"05721383",
  1440 => x"712b7208",
  1441 => x"07720c53",
  1442 => x"53800b80",
  1443 => x"dfb80c80",
  1444 => x"0b80dfb4",
  1445 => x"0c80e2f4",
  1446 => x"51afd62d",
  1447 => x"80e18008",
  1448 => x"ff24feea",
  1449 => x"38aae62d",
  1450 => x"80e18008",
  1451 => x"802e81b0",
  1452 => x"38815980",
  1453 => x"0b80dfb0",
  1454 => x"0880dfac",
  1455 => x"0880dee0",
  1456 => x"5a5c5c58",
  1457 => x"7a79067a",
  1458 => x"7a065452",
  1459 => x"71732e80",
  1460 => x"f8387209",
  1461 => x"81057074",
  1462 => x"07802580",
  1463 => x"decc1a80",
  1464 => x"f52d7084",
  1465 => x"2c718f06",
  1466 => x"58535757",
  1467 => x"5275802e",
  1468 => x"a3387184",
  1469 => x"2980de8c",
  1470 => x"05741583",
  1471 => x"712b7208",
  1472 => x"07720c54",
  1473 => x"527680e0",
  1474 => x"2d810552",
  1475 => x"7177818a",
  1476 => x"2daeaa04",
  1477 => x"71842980",
  1478 => x"de8c0574",
  1479 => x"1581712b",
  1480 => x"70097308",
  1481 => x"06730c51",
  1482 => x"53537485",
  1483 => x"32700981",
  1484 => x"05708025",
  1485 => x"51515275",
  1486 => x"802e8e38",
  1487 => x"81707306",
  1488 => x"53537180",
  1489 => x"2e833872",
  1490 => x"5c781081",
  1491 => x"19821959",
  1492 => x"59599078",
  1493 => x"25feed38",
  1494 => x"80dfac08",
  1495 => x"80dfb00c",
  1496 => x"7b80e180",
  1497 => x"0c02b005",
  1498 => x"0d0402f8",
  1499 => x"050d80de",
  1500 => x"8c528f51",
  1501 => x"80727084",
  1502 => x"05540cff",
  1503 => x"11517080",
  1504 => x"25f23802",
  1505 => x"88050d04",
  1506 => x"02f0050d",
  1507 => x"7551aae0",
  1508 => x"2d70822c",
  1509 => x"fc0680de",
  1510 => x"8c117210",
  1511 => x"9e067108",
  1512 => x"70722a70",
  1513 => x"83068274",
  1514 => x"2b700974",
  1515 => x"06760c54",
  1516 => x"51565753",
  1517 => x"5153aada",
  1518 => x"2d7180e1",
  1519 => x"800c0290",
  1520 => x"050d0402",
  1521 => x"fc050d72",
  1522 => x"5180710c",
  1523 => x"800b8412",
  1524 => x"0c028405",
  1525 => x"0d0402f0",
  1526 => x"050d7570",
  1527 => x"08841208",
  1528 => x"535353ff",
  1529 => x"5471712e",
  1530 => x"a838aae0",
  1531 => x"2d841308",
  1532 => x"70842914",
  1533 => x"88117008",
  1534 => x"7081ff06",
  1535 => x"84180881",
  1536 => x"11870684",
  1537 => x"1a0c5351",
  1538 => x"55515151",
  1539 => x"aada2d71",
  1540 => x"547380e1",
  1541 => x"800c0290",
  1542 => x"050d0402",
  1543 => x"f8050daa",
  1544 => x"e02de008",
  1545 => x"708b2a70",
  1546 => x"81065152",
  1547 => x"5270802e",
  1548 => x"a13880e2",
  1549 => x"f4087084",
  1550 => x"2980e2fc",
  1551 => x"057381ff",
  1552 => x"06710c51",
  1553 => x"5180e2f4",
  1554 => x"08811187",
  1555 => x"0680e2f4",
  1556 => x"0c51800b",
  1557 => x"80e39c0c",
  1558 => x"aad22daa",
  1559 => x"da2d0288",
  1560 => x"050d0402",
  1561 => x"fc050daa",
  1562 => x"e02d810b",
  1563 => x"80e39c0c",
  1564 => x"aada2d80",
  1565 => x"e39c0851",
  1566 => x"70f93802",
  1567 => x"84050d04",
  1568 => x"02fc050d",
  1569 => x"80e2f451",
  1570 => x"afc32dae",
  1571 => x"ea2db09b",
  1572 => x"51aace2d",
  1573 => x"0284050d",
  1574 => x"0480e3a8",
  1575 => x"0880e180",
  1576 => x"0c0402fc",
  1577 => x"050d810b",
  1578 => x"80dfc00c",
  1579 => x"8151858d",
  1580 => x"2d028405",
  1581 => x"0d0402fc",
  1582 => x"050db1c0",
  1583 => x"04ac852d",
  1584 => x"80f651af",
  1585 => x"882d80e1",
  1586 => x"8008f238",
  1587 => x"80da51af",
  1588 => x"882d80e1",
  1589 => x"8008e638",
  1590 => x"80e18008",
  1591 => x"80dfc00c",
  1592 => x"80e18008",
  1593 => x"51858d2d",
  1594 => x"0284050d",
  1595 => x"0402ec05",
  1596 => x"0d765480",
  1597 => x"52870b88",
  1598 => x"1580f52d",
  1599 => x"56537472",
  1600 => x"248338a0",
  1601 => x"53725183",
  1602 => x"842d8112",
  1603 => x"8b1580f5",
  1604 => x"2d545272",
  1605 => x"7225de38",
  1606 => x"0294050d",
  1607 => x"0402f005",
  1608 => x"0d80e3a8",
  1609 => x"085481f9",
  1610 => x"2d800b80",
  1611 => x"e3ac0c73",
  1612 => x"08802e81",
  1613 => x"8938820b",
  1614 => x"80e1940c",
  1615 => x"80e3ac08",
  1616 => x"8f0680e1",
  1617 => x"900c7308",
  1618 => x"5271832e",
  1619 => x"96387183",
  1620 => x"26893871",
  1621 => x"812eb038",
  1622 => x"b3a70471",
  1623 => x"852ea038",
  1624 => x"b3a70488",
  1625 => x"1480f52d",
  1626 => x"84150880",
  1627 => x"dae45354",
  1628 => x"5286a02d",
  1629 => x"71842913",
  1630 => x"70085252",
  1631 => x"b3ab0473",
  1632 => x"51b1ed2d",
  1633 => x"b3a70480",
  1634 => x"dfbc0888",
  1635 => x"15082c70",
  1636 => x"81065152",
  1637 => x"71802e88",
  1638 => x"3880dae8",
  1639 => x"51b3a404",
  1640 => x"80daec51",
  1641 => x"86a02d84",
  1642 => x"14085186",
  1643 => x"a02d80e3",
  1644 => x"ac088105",
  1645 => x"80e3ac0c",
  1646 => x"8c1454b2",
  1647 => x"af040290",
  1648 => x"050d0471",
  1649 => x"80e3a80c",
  1650 => x"b29d2d80",
  1651 => x"e3ac08ff",
  1652 => x"0580e3b0",
  1653 => x"0c0402e8",
  1654 => x"050d80e3",
  1655 => x"a80880e3",
  1656 => x"b4085755",
  1657 => x"80f651af",
  1658 => x"882d80e1",
  1659 => x"8008812a",
  1660 => x"70810651",
  1661 => x"5271802e",
  1662 => x"a438b480",
  1663 => x"04ac852d",
  1664 => x"80f651af",
  1665 => x"882d80e1",
  1666 => x"8008f238",
  1667 => x"80dfc008",
  1668 => x"81327080",
  1669 => x"dfc00c70",
  1670 => x"5252858d",
  1671 => x"2d800b80",
  1672 => x"e3a00c80",
  1673 => x"0b80e3a4",
  1674 => x"0c80dfc0",
  1675 => x"08838d38",
  1676 => x"80da51af",
  1677 => x"882d80e1",
  1678 => x"8008802e",
  1679 => x"8c3880e3",
  1680 => x"a0088180",
  1681 => x"0780e3a0",
  1682 => x"0c80d951",
  1683 => x"af882d80",
  1684 => x"e1800880",
  1685 => x"2e8c3880",
  1686 => x"e3a00880",
  1687 => x"c00780e3",
  1688 => x"a00c8194",
  1689 => x"51af882d",
  1690 => x"80e18008",
  1691 => x"802e8b38",
  1692 => x"80e3a008",
  1693 => x"900780e3",
  1694 => x"a00c8191",
  1695 => x"51af882d",
  1696 => x"80e18008",
  1697 => x"802e8b38",
  1698 => x"80e3a008",
  1699 => x"a00780e3",
  1700 => x"a00c81f5",
  1701 => x"51af882d",
  1702 => x"80e18008",
  1703 => x"802e8b38",
  1704 => x"80e3a008",
  1705 => x"810780e3",
  1706 => x"a00c81f2",
  1707 => x"51af882d",
  1708 => x"80e18008",
  1709 => x"802e8b38",
  1710 => x"80e3a008",
  1711 => x"820780e3",
  1712 => x"a00c81eb",
  1713 => x"51af882d",
  1714 => x"80e18008",
  1715 => x"802e8b38",
  1716 => x"80e3a008",
  1717 => x"840780e3",
  1718 => x"a00c81f4",
  1719 => x"51af882d",
  1720 => x"80e18008",
  1721 => x"802e8b38",
  1722 => x"80e3a008",
  1723 => x"880780e3",
  1724 => x"a00c80d8",
  1725 => x"51af882d",
  1726 => x"80e18008",
  1727 => x"802e8c38",
  1728 => x"80e3a408",
  1729 => x"81800780",
  1730 => x"e3a40c92",
  1731 => x"51af882d",
  1732 => x"80e18008",
  1733 => x"802e8c38",
  1734 => x"80e3a408",
  1735 => x"80c00780",
  1736 => x"e3a40c94",
  1737 => x"51af882d",
  1738 => x"80e18008",
  1739 => x"802e8b38",
  1740 => x"80e3a408",
  1741 => x"900780e3",
  1742 => x"a40c9151",
  1743 => x"af882d80",
  1744 => x"e1800880",
  1745 => x"2e8b3880",
  1746 => x"e3a408a0",
  1747 => x"0780e3a4",
  1748 => x"0c9d51af",
  1749 => x"882d80e1",
  1750 => x"8008802e",
  1751 => x"8b3880e3",
  1752 => x"a4088107",
  1753 => x"80e3a40c",
  1754 => x"9b51af88",
  1755 => x"2d80e180",
  1756 => x"08802e8b",
  1757 => x"3880e3a4",
  1758 => x"08820780",
  1759 => x"e3a40c9c",
  1760 => x"51af882d",
  1761 => x"80e18008",
  1762 => x"802e8b38",
  1763 => x"80e3a408",
  1764 => x"840780e3",
  1765 => x"a40ca351",
  1766 => x"af882d80",
  1767 => x"e1800880",
  1768 => x"2e8b3880",
  1769 => x"e3a40888",
  1770 => x"0780e3a4",
  1771 => x"0c81fd51",
  1772 => x"af882d81",
  1773 => x"fa51af88",
  1774 => x"2dbd9104",
  1775 => x"81f551af",
  1776 => x"882d80e1",
  1777 => x"8008812a",
  1778 => x"70810651",
  1779 => x"5271802e",
  1780 => x"b33880e3",
  1781 => x"b0085271",
  1782 => x"802e8a38",
  1783 => x"ff1280e3",
  1784 => x"b00cb884",
  1785 => x"0480e3ac",
  1786 => x"081080e3",
  1787 => x"ac080570",
  1788 => x"84291651",
  1789 => x"52881208",
  1790 => x"802e8938",
  1791 => x"ff518812",
  1792 => x"0852712d",
  1793 => x"81f251af",
  1794 => x"882d80e1",
  1795 => x"8008812a",
  1796 => x"70810651",
  1797 => x"5271802e",
  1798 => x"b43880e3",
  1799 => x"ac08ff11",
  1800 => x"80e3b008",
  1801 => x"56535373",
  1802 => x"72258a38",
  1803 => x"811480e3",
  1804 => x"b00cb8cd",
  1805 => x"04721013",
  1806 => x"70842916",
  1807 => x"51528812",
  1808 => x"08802e89",
  1809 => x"38fe5188",
  1810 => x"12085271",
  1811 => x"2d81fd51",
  1812 => x"af882d80",
  1813 => x"e1800881",
  1814 => x"2a708106",
  1815 => x"51527180",
  1816 => x"2eb13880",
  1817 => x"e3b00880",
  1818 => x"2e8a3880",
  1819 => x"0b80e3b0",
  1820 => x"0cb99304",
  1821 => x"80e3ac08",
  1822 => x"1080e3ac",
  1823 => x"08057084",
  1824 => x"29165152",
  1825 => x"88120880",
  1826 => x"2e8938fd",
  1827 => x"51881208",
  1828 => x"52712d81",
  1829 => x"fa51af88",
  1830 => x"2d80e180",
  1831 => x"08812a70",
  1832 => x"81065152",
  1833 => x"71802eb1",
  1834 => x"3880e3ac",
  1835 => x"08ff1154",
  1836 => x"5280e3b0",
  1837 => x"08732589",
  1838 => x"387280e3",
  1839 => x"b00cb9d9",
  1840 => x"04711012",
  1841 => x"70842916",
  1842 => x"51528812",
  1843 => x"08802e89",
  1844 => x"38fc5188",
  1845 => x"12085271",
  1846 => x"2d80e3b0",
  1847 => x"08705354",
  1848 => x"73802e8a",
  1849 => x"388c15ff",
  1850 => x"155555b9",
  1851 => x"e004820b",
  1852 => x"80e1940c",
  1853 => x"718f0680",
  1854 => x"e1900c81",
  1855 => x"eb51af88",
  1856 => x"2d80e180",
  1857 => x"08812a70",
  1858 => x"81065152",
  1859 => x"71802ead",
  1860 => x"38740885",
  1861 => x"2e098106",
  1862 => x"a4388815",
  1863 => x"80f52dff",
  1864 => x"05527188",
  1865 => x"1681b72d",
  1866 => x"71982b52",
  1867 => x"71802588",
  1868 => x"38800b88",
  1869 => x"1681b72d",
  1870 => x"7451b1ed",
  1871 => x"2d81f451",
  1872 => x"af882d80",
  1873 => x"e1800881",
  1874 => x"2a708106",
  1875 => x"51527180",
  1876 => x"2eb33874",
  1877 => x"08852e09",
  1878 => x"8106aa38",
  1879 => x"881580f5",
  1880 => x"2d810552",
  1881 => x"71881681",
  1882 => x"b72d7181",
  1883 => x"ff068b16",
  1884 => x"80f52d54",
  1885 => x"52727227",
  1886 => x"87387288",
  1887 => x"1681b72d",
  1888 => x"7451b1ed",
  1889 => x"2d80da51",
  1890 => x"af882d80",
  1891 => x"e1800881",
  1892 => x"2a708106",
  1893 => x"51527180",
  1894 => x"2e81ad38",
  1895 => x"80e3a808",
  1896 => x"80e3b008",
  1897 => x"55537380",
  1898 => x"2e8a388c",
  1899 => x"13ff1555",
  1900 => x"53bba604",
  1901 => x"72085271",
  1902 => x"822ea638",
  1903 => x"71822689",
  1904 => x"3871812e",
  1905 => x"aa38bcc8",
  1906 => x"0471832e",
  1907 => x"b4387184",
  1908 => x"2e098106",
  1909 => x"80f23888",
  1910 => x"130851b3",
  1911 => x"c32dbcc8",
  1912 => x"0480e3b0",
  1913 => x"08518813",
  1914 => x"0852712d",
  1915 => x"bcc80481",
  1916 => x"0b881408",
  1917 => x"2b80dfbc",
  1918 => x"083280df",
  1919 => x"bc0cbc9c",
  1920 => x"04881380",
  1921 => x"f52d8105",
  1922 => x"8b1480f5",
  1923 => x"2d535471",
  1924 => x"74248338",
  1925 => x"80547388",
  1926 => x"1481b72d",
  1927 => x"b29d2dbc",
  1928 => x"c8047508",
  1929 => x"802ea438",
  1930 => x"750851af",
  1931 => x"882d80e1",
  1932 => x"80088106",
  1933 => x"5271802e",
  1934 => x"8c3880e3",
  1935 => x"b0085184",
  1936 => x"16085271",
  1937 => x"2d881656",
  1938 => x"75d83880",
  1939 => x"54800b80",
  1940 => x"e1940c73",
  1941 => x"8f0680e1",
  1942 => x"900ca052",
  1943 => x"7380e3b0",
  1944 => x"082e0981",
  1945 => x"06993880",
  1946 => x"e3ac08ff",
  1947 => x"05743270",
  1948 => x"09810570",
  1949 => x"72079f2a",
  1950 => x"91713151",
  1951 => x"51535371",
  1952 => x"5183842d",
  1953 => x"8114548e",
  1954 => x"7425c238",
  1955 => x"80dfc008",
  1956 => x"527180e1",
  1957 => x"800c0298",
  1958 => x"050d0402",
  1959 => x"f4050dd4",
  1960 => x"5281ff72",
  1961 => x"0c710853",
  1962 => x"81ff720c",
  1963 => x"72882b83",
  1964 => x"fe800672",
  1965 => x"087081ff",
  1966 => x"06515253",
  1967 => x"81ff720c",
  1968 => x"72710788",
  1969 => x"2b720870",
  1970 => x"81ff0651",
  1971 => x"525381ff",
  1972 => x"720c7271",
  1973 => x"07882b72",
  1974 => x"087081ff",
  1975 => x"06720780",
  1976 => x"e1800c52",
  1977 => x"53028c05",
  1978 => x"0d0402f4",
  1979 => x"050d7476",
  1980 => x"7181ff06",
  1981 => x"d40c5353",
  1982 => x"80e3b808",
  1983 => x"85387189",
  1984 => x"2b527198",
  1985 => x"2ad40c71",
  1986 => x"902a7081",
  1987 => x"ff06d40c",
  1988 => x"5171882a",
  1989 => x"7081ff06",
  1990 => x"d40c5171",
  1991 => x"81ff06d4",
  1992 => x"0c72902a",
  1993 => x"7081ff06",
  1994 => x"d40c51d4",
  1995 => x"087081ff",
  1996 => x"06515182",
  1997 => x"b8bf5270",
  1998 => x"81ff2e09",
  1999 => x"81069438",
  2000 => x"81ff0bd4",
  2001 => x"0cd40870",
  2002 => x"81ff06ff",
  2003 => x"14545151",
  2004 => x"71e53870",
  2005 => x"80e1800c",
  2006 => x"028c050d",
  2007 => x"0402fc05",
  2008 => x"0d81c751",
  2009 => x"81ff0bd4",
  2010 => x"0cff1151",
  2011 => x"708025f4",
  2012 => x"38028405",
  2013 => x"0d0402f4",
  2014 => x"050d81ff",
  2015 => x"0bd40c93",
  2016 => x"53805287",
  2017 => x"fc80c151",
  2018 => x"bdea2d80",
  2019 => x"e180088b",
  2020 => x"3881ff0b",
  2021 => x"d40c8153",
  2022 => x"bfa404be",
  2023 => x"dd2dff13",
  2024 => x"5372de38",
  2025 => x"7280e180",
  2026 => x"0c028c05",
  2027 => x"0d0402ec",
  2028 => x"050d810b",
  2029 => x"80e3b80c",
  2030 => x"8454d008",
  2031 => x"708f2a70",
  2032 => x"81065151",
  2033 => x"5372f338",
  2034 => x"72d00cbe",
  2035 => x"dd2d80da",
  2036 => x"f05186a0",
  2037 => x"2dd00870",
  2038 => x"8f2a7081",
  2039 => x"06515153",
  2040 => x"72f33881",
  2041 => x"0bd00cb1",
  2042 => x"53805284",
  2043 => x"d480c051",
  2044 => x"bdea2d80",
  2045 => x"e1800881",
  2046 => x"2e943872",
  2047 => x"822e80c0",
  2048 => x"38ff1353",
  2049 => x"72e338ff",
  2050 => x"145473ff",
  2051 => x"ad38bedd",
  2052 => x"2d83aa52",
  2053 => x"849c80c8",
  2054 => x"51bdea2d",
  2055 => x"80e18008",
  2056 => x"812e0981",
  2057 => x"069338bd",
  2058 => x"9b2d80e1",
  2059 => x"800883ff",
  2060 => x"ff065372",
  2061 => x"83aa2ea2",
  2062 => x"38bef62d",
  2063 => x"80c0d404",
  2064 => x"80dafc51",
  2065 => x"86a02d80",
  2066 => x"5380c2ac",
  2067 => x"0480db94",
  2068 => x"5186a02d",
  2069 => x"805480c1",
  2070 => x"fd0481ff",
  2071 => x"0bd40cb1",
  2072 => x"54bedd2d",
  2073 => x"8fcf5380",
  2074 => x"5287fc80",
  2075 => x"f751bdea",
  2076 => x"2d80e180",
  2077 => x"085580e1",
  2078 => x"8008812e",
  2079 => x"0981069c",
  2080 => x"3881ff0b",
  2081 => x"d40c820a",
  2082 => x"52849c80",
  2083 => x"e951bdea",
  2084 => x"2d80e180",
  2085 => x"08802e8e",
  2086 => x"38bedd2d",
  2087 => x"ff135372",
  2088 => x"c63880c1",
  2089 => x"f00481ff",
  2090 => x"0bd40c80",
  2091 => x"e1800852",
  2092 => x"87fc80fa",
  2093 => x"51bdea2d",
  2094 => x"80e18008",
  2095 => x"b33881ff",
  2096 => x"0bd40cd4",
  2097 => x"085381ff",
  2098 => x"0bd40c81",
  2099 => x"ff0bd40c",
  2100 => x"81ff0bd4",
  2101 => x"0c81ff0b",
  2102 => x"d40c7286",
  2103 => x"2a708106",
  2104 => x"76565153",
  2105 => x"72973880",
  2106 => x"e1800854",
  2107 => x"80c1fd04",
  2108 => x"73822efe",
  2109 => x"d838ff14",
  2110 => x"5473fee5",
  2111 => x"387380e3",
  2112 => x"b80c738b",
  2113 => x"38815287",
  2114 => x"fc80d051",
  2115 => x"bdea2d81",
  2116 => x"ff0bd40c",
  2117 => x"d008708f",
  2118 => x"2a708106",
  2119 => x"51515372",
  2120 => x"f33872d0",
  2121 => x"0c81ff0b",
  2122 => x"d40c8153",
  2123 => x"7280e180",
  2124 => x"0c029405",
  2125 => x"0d0402e8",
  2126 => x"050d7855",
  2127 => x"805681ff",
  2128 => x"0bd40cd0",
  2129 => x"08708f2a",
  2130 => x"70810651",
  2131 => x"515372f3",
  2132 => x"3882810b",
  2133 => x"d00c81ff",
  2134 => x"0bd40c77",
  2135 => x"5287fc80",
  2136 => x"d151bdea",
  2137 => x"2d80dbc6",
  2138 => x"df5480e1",
  2139 => x"8008802e",
  2140 => x"8c3880db",
  2141 => x"b45186a0",
  2142 => x"2d80c3d2",
  2143 => x"0481ff0b",
  2144 => x"d40cd408",
  2145 => x"7081ff06",
  2146 => x"51537281",
  2147 => x"fe2e0981",
  2148 => x"069f3880",
  2149 => x"ff53bd9b",
  2150 => x"2d80e180",
  2151 => x"08757084",
  2152 => x"05570cff",
  2153 => x"13537280",
  2154 => x"25ec3881",
  2155 => x"5680c3b7",
  2156 => x"04ff1454",
  2157 => x"73c73881",
  2158 => x"ff0bd40c",
  2159 => x"81ff0bd4",
  2160 => x"0cd00870",
  2161 => x"8f2a7081",
  2162 => x"06515153",
  2163 => x"72f33872",
  2164 => x"d00c7580",
  2165 => x"e1800c02",
  2166 => x"98050d04",
  2167 => x"02e8050d",
  2168 => x"77797b58",
  2169 => x"55558053",
  2170 => x"727625a5",
  2171 => x"38747081",
  2172 => x"055680f5",
  2173 => x"2d747081",
  2174 => x"055680f5",
  2175 => x"2d525271",
  2176 => x"712e8738",
  2177 => x"815180c4",
  2178 => x"93048113",
  2179 => x"5380c3e8",
  2180 => x"04805170",
  2181 => x"80e1800c",
  2182 => x"0298050d",
  2183 => x"0402ec05",
  2184 => x"0d765574",
  2185 => x"802e80c4",
  2186 => x"389a1580",
  2187 => x"e02d5180",
  2188 => x"d2d72d80",
  2189 => x"e1800880",
  2190 => x"e1800880",
  2191 => x"e9ec0c80",
  2192 => x"e1800854",
  2193 => x"5480e9c8",
  2194 => x"08802e9b",
  2195 => x"38941580",
  2196 => x"e02d5180",
  2197 => x"d2d72d80",
  2198 => x"e1800890",
  2199 => x"2b83fff0",
  2200 => x"0a067075",
  2201 => x"07515372",
  2202 => x"80e9ec0c",
  2203 => x"80e9ec08",
  2204 => x"5372802e",
  2205 => x"9e3880e9",
  2206 => x"c008fe14",
  2207 => x"712980e9",
  2208 => x"d4080580",
  2209 => x"e9f00c70",
  2210 => x"842b80e9",
  2211 => x"cc0c5480",
  2212 => x"c5c20480",
  2213 => x"e9d80880",
  2214 => x"e9ec0c80",
  2215 => x"e9dc0880",
  2216 => x"e9f00c80",
  2217 => x"e9c80880",
  2218 => x"2e8c3880",
  2219 => x"e9c00884",
  2220 => x"2b5380c5",
  2221 => x"bd0480e9",
  2222 => x"e008842b",
  2223 => x"537280e9",
  2224 => x"cc0c0294",
  2225 => x"050d0402",
  2226 => x"d8050d80",
  2227 => x"0b80e9c8",
  2228 => x"0c8454bf",
  2229 => x"ae2d80e1",
  2230 => x"8008802e",
  2231 => x"993880e3",
  2232 => x"bc528051",
  2233 => x"80c2b62d",
  2234 => x"80e18008",
  2235 => x"802e8738",
  2236 => x"fe5480c5",
  2237 => x"fe04ff14",
  2238 => x"54738024",
  2239 => x"d638738e",
  2240 => x"3880dbc4",
  2241 => x"5186a02d",
  2242 => x"735580cb",
  2243 => x"e2048056",
  2244 => x"810b80e9",
  2245 => x"f40c8853",
  2246 => x"80dbd852",
  2247 => x"80e3f251",
  2248 => x"80c3dc2d",
  2249 => x"80e18008",
  2250 => x"762e0981",
  2251 => x"06893880",
  2252 => x"e1800880",
  2253 => x"e9f40c88",
  2254 => x"5380dbe4",
  2255 => x"5280e48e",
  2256 => x"5180c3dc",
  2257 => x"2d80e180",
  2258 => x"08893880",
  2259 => x"e1800880",
  2260 => x"e9f40c80",
  2261 => x"e9f40880",
  2262 => x"2e818538",
  2263 => x"80e7820b",
  2264 => x"80f52d80",
  2265 => x"e7830b80",
  2266 => x"f52d7198",
  2267 => x"2b71902b",
  2268 => x"0780e784",
  2269 => x"0b80f52d",
  2270 => x"70882b72",
  2271 => x"0780e785",
  2272 => x"0b80f52d",
  2273 => x"710780e7",
  2274 => x"ba0b80f5",
  2275 => x"2d80e7bb",
  2276 => x"0b80f52d",
  2277 => x"71882b07",
  2278 => x"535f5452",
  2279 => x"5a565755",
  2280 => x"7381abaa",
  2281 => x"2e098106",
  2282 => x"90387551",
  2283 => x"80d2a62d",
  2284 => x"80e18008",
  2285 => x"5680c7c8",
  2286 => x"047382d4",
  2287 => x"d52e8938",
  2288 => x"80dbf051",
  2289 => x"80c89804",
  2290 => x"80e3bc52",
  2291 => x"755180c2",
  2292 => x"b62d80e1",
  2293 => x"80085580",
  2294 => x"e1800880",
  2295 => x"2e848338",
  2296 => x"885380db",
  2297 => x"e45280e4",
  2298 => x"8e5180c3",
  2299 => x"dc2d80e1",
  2300 => x"80088b38",
  2301 => x"810b80e9",
  2302 => x"c80c80c8",
  2303 => x"9f048853",
  2304 => x"80dbd852",
  2305 => x"80e3f251",
  2306 => x"80c3dc2d",
  2307 => x"80e18008",
  2308 => x"802e8c38",
  2309 => x"80dc8451",
  2310 => x"86a02d80",
  2311 => x"c8fe0480",
  2312 => x"e7ba0b80",
  2313 => x"f52d5473",
  2314 => x"80d52e09",
  2315 => x"810680ce",
  2316 => x"3880e7bb",
  2317 => x"0b80f52d",
  2318 => x"547381aa",
  2319 => x"2e098106",
  2320 => x"bd38800b",
  2321 => x"80e3bc0b",
  2322 => x"80f52d56",
  2323 => x"547481e9",
  2324 => x"2e833881",
  2325 => x"547481eb",
  2326 => x"2e8c3880",
  2327 => x"5573752e",
  2328 => x"09810682",
  2329 => x"fd3880e3",
  2330 => x"c70b80f5",
  2331 => x"2d55748e",
  2332 => x"3880e3c8",
  2333 => x"0b80f52d",
  2334 => x"5473822e",
  2335 => x"87388055",
  2336 => x"80cbe204",
  2337 => x"80e3c90b",
  2338 => x"80f52d70",
  2339 => x"80e9c00c",
  2340 => x"ff0580e9",
  2341 => x"c40c80e3",
  2342 => x"ca0b80f5",
  2343 => x"2d80e3cb",
  2344 => x"0b80f52d",
  2345 => x"58760577",
  2346 => x"82802905",
  2347 => x"7080e9d0",
  2348 => x"0c80e3cc",
  2349 => x"0b80f52d",
  2350 => x"7080e9e4",
  2351 => x"0c80e9c8",
  2352 => x"08595758",
  2353 => x"76802e81",
  2354 => x"b9388853",
  2355 => x"80dbe452",
  2356 => x"80e48e51",
  2357 => x"80c3dc2d",
  2358 => x"80e18008",
  2359 => x"82843880",
  2360 => x"e9c00870",
  2361 => x"842b80e9",
  2362 => x"cc0c7080",
  2363 => x"e9e00c80",
  2364 => x"e3e10b80",
  2365 => x"f52d80e3",
  2366 => x"e00b80f5",
  2367 => x"2d718280",
  2368 => x"290580e3",
  2369 => x"e20b80f5",
  2370 => x"2d708480",
  2371 => x"80291280",
  2372 => x"e3e30b80",
  2373 => x"f52d7081",
  2374 => x"800a2912",
  2375 => x"7080e9e8",
  2376 => x"0c80e9e4",
  2377 => x"08712980",
  2378 => x"e9d00805",
  2379 => x"7080e9d4",
  2380 => x"0c80e3e9",
  2381 => x"0b80f52d",
  2382 => x"80e3e80b",
  2383 => x"80f52d71",
  2384 => x"82802905",
  2385 => x"80e3ea0b",
  2386 => x"80f52d70",
  2387 => x"84808029",
  2388 => x"1280e3eb",
  2389 => x"0b80f52d",
  2390 => x"70982b81",
  2391 => x"f00a0672",
  2392 => x"057080e9",
  2393 => x"d80cfe11",
  2394 => x"7e297705",
  2395 => x"80e9dc0c",
  2396 => x"52595243",
  2397 => x"545e5152",
  2398 => x"59525d57",
  2399 => x"595780cb",
  2400 => x"da0480e3",
  2401 => x"ce0b80f5",
  2402 => x"2d80e3cd",
  2403 => x"0b80f52d",
  2404 => x"71828029",
  2405 => x"057080e9",
  2406 => x"cc0c70a0",
  2407 => x"2983ff05",
  2408 => x"70892a70",
  2409 => x"80e9e00c",
  2410 => x"80e3d30b",
  2411 => x"80f52d80",
  2412 => x"e3d20b80",
  2413 => x"f52d7182",
  2414 => x"80290570",
  2415 => x"80e9e80c",
  2416 => x"7b71291e",
  2417 => x"7080e9dc",
  2418 => x"0c7d80e9",
  2419 => x"d80c7305",
  2420 => x"80e9d40c",
  2421 => x"555e5151",
  2422 => x"55558051",
  2423 => x"80c49d2d",
  2424 => x"81557480",
  2425 => x"e1800c02",
  2426 => x"a8050d04",
  2427 => x"02ec050d",
  2428 => x"7670872c",
  2429 => x"7180ff06",
  2430 => x"55565480",
  2431 => x"e9c8088a",
  2432 => x"3873882c",
  2433 => x"7481ff06",
  2434 => x"545580e3",
  2435 => x"bc5280e9",
  2436 => x"d0081551",
  2437 => x"80c2b62d",
  2438 => x"80e18008",
  2439 => x"5480e180",
  2440 => x"08802ebb",
  2441 => x"3880e9c8",
  2442 => x"08802e9c",
  2443 => x"38728429",
  2444 => x"80e3bc05",
  2445 => x"70085253",
  2446 => x"80d2a62d",
  2447 => x"80e18008",
  2448 => x"f00a0653",
  2449 => x"80ccdd04",
  2450 => x"721080e3",
  2451 => x"bc057080",
  2452 => x"e02d5253",
  2453 => x"80d2d72d",
  2454 => x"80e18008",
  2455 => x"53725473",
  2456 => x"80e1800c",
  2457 => x"0294050d",
  2458 => x"0402e005",
  2459 => x"0d797084",
  2460 => x"2c80e9f0",
  2461 => x"0805718f",
  2462 => x"06525553",
  2463 => x"728b3880",
  2464 => x"e3bc5273",
  2465 => x"5180c2b6",
  2466 => x"2d72a029",
  2467 => x"80e3bc05",
  2468 => x"54807480",
  2469 => x"f52d5653",
  2470 => x"74732e83",
  2471 => x"38815374",
  2472 => x"81e52e81",
  2473 => x"f5388170",
  2474 => x"74065458",
  2475 => x"72802e81",
  2476 => x"e9388b14",
  2477 => x"80f52d70",
  2478 => x"832a7906",
  2479 => x"5856769c",
  2480 => x"3880dfc4",
  2481 => x"08537289",
  2482 => x"387280e7",
  2483 => x"bc0b81b7",
  2484 => x"2d7680df",
  2485 => x"c40c7353",
  2486 => x"80cf9c04",
  2487 => x"758f2e09",
  2488 => x"810681b6",
  2489 => x"38749f06",
  2490 => x"8d2980e7",
  2491 => x"af115153",
  2492 => x"811480f5",
  2493 => x"2d737081",
  2494 => x"055581b7",
  2495 => x"2d831480",
  2496 => x"f52d7370",
  2497 => x"81055581",
  2498 => x"b72d8514",
  2499 => x"80f52d73",
  2500 => x"70810555",
  2501 => x"81b72d87",
  2502 => x"1480f52d",
  2503 => x"73708105",
  2504 => x"5581b72d",
  2505 => x"891480f5",
  2506 => x"2d737081",
  2507 => x"055581b7",
  2508 => x"2d8e1480",
  2509 => x"f52d7370",
  2510 => x"81055581",
  2511 => x"b72d9014",
  2512 => x"80f52d73",
  2513 => x"70810555",
  2514 => x"81b72d92",
  2515 => x"1480f52d",
  2516 => x"73708105",
  2517 => x"5581b72d",
  2518 => x"941480f5",
  2519 => x"2d737081",
  2520 => x"055581b7",
  2521 => x"2d961480",
  2522 => x"f52d7370",
  2523 => x"81055581",
  2524 => x"b72d9814",
  2525 => x"80f52d73",
  2526 => x"70810555",
  2527 => x"81b72d9c",
  2528 => x"1480f52d",
  2529 => x"73708105",
  2530 => x"5581b72d",
  2531 => x"9e1480f5",
  2532 => x"2d7381b7",
  2533 => x"2d7780df",
  2534 => x"c40c8053",
  2535 => x"7280e180",
  2536 => x"0c02a005",
  2537 => x"0d0402cc",
  2538 => x"050d7e60",
  2539 => x"5e5a800b",
  2540 => x"80e9ec08",
  2541 => x"80e9f008",
  2542 => x"595c5680",
  2543 => x"5880e9cc",
  2544 => x"08782e81",
  2545 => x"be38778f",
  2546 => x"06a01757",
  2547 => x"54739238",
  2548 => x"80e3bc52",
  2549 => x"76518117",
  2550 => x"5780c2b6",
  2551 => x"2d80e3bc",
  2552 => x"56807680",
  2553 => x"f52d5654",
  2554 => x"74742e83",
  2555 => x"38815474",
  2556 => x"81e52e81",
  2557 => x"82388170",
  2558 => x"7506555c",
  2559 => x"73802e80",
  2560 => x"f6388b16",
  2561 => x"80f52d98",
  2562 => x"06597880",
  2563 => x"ea388b53",
  2564 => x"7c527551",
  2565 => x"80c3dc2d",
  2566 => x"80e18008",
  2567 => x"80d9389c",
  2568 => x"16085180",
  2569 => x"d2a62d80",
  2570 => x"e1800884",
  2571 => x"1b0c9a16",
  2572 => x"80e02d51",
  2573 => x"80d2d72d",
  2574 => x"80e18008",
  2575 => x"80e18008",
  2576 => x"881c0c80",
  2577 => x"e1800855",
  2578 => x"5580e9c8",
  2579 => x"08802e9a",
  2580 => x"38941680",
  2581 => x"e02d5180",
  2582 => x"d2d72d80",
  2583 => x"e1800890",
  2584 => x"2b83fff0",
  2585 => x"0a067016",
  2586 => x"51547388",
  2587 => x"1b0c787a",
  2588 => x"0c7b5480",
  2589 => x"d1c10481",
  2590 => x"185880e9",
  2591 => x"cc087826",
  2592 => x"fec43880",
  2593 => x"e9c80880",
  2594 => x"2eb5387a",
  2595 => x"5180cbec",
  2596 => x"2d80e180",
  2597 => x"0880e180",
  2598 => x"0880ffff",
  2599 => x"fff80655",
  2600 => x"5b7380ff",
  2601 => x"fffff82e",
  2602 => x"963880e1",
  2603 => x"8008fe05",
  2604 => x"80e9c008",
  2605 => x"2980e9d4",
  2606 => x"08055780",
  2607 => x"cfbb0480",
  2608 => x"547380e1",
  2609 => x"800c02b4",
  2610 => x"050d0402",
  2611 => x"f4050d74",
  2612 => x"70088105",
  2613 => x"710c7008",
  2614 => x"80e9c408",
  2615 => x"06535371",
  2616 => x"90388813",
  2617 => x"085180cb",
  2618 => x"ec2d80e1",
  2619 => x"80088814",
  2620 => x"0c810b80",
  2621 => x"e1800c02",
  2622 => x"8c050d04",
  2623 => x"02f0050d",
  2624 => x"75881108",
  2625 => x"fe0580e9",
  2626 => x"c0082980",
  2627 => x"e9d40811",
  2628 => x"720880e9",
  2629 => x"c4080605",
  2630 => x"79555354",
  2631 => x"5480c2b6",
  2632 => x"2d029005",
  2633 => x"0d0402f4",
  2634 => x"050d7470",
  2635 => x"882a83fe",
  2636 => x"80067072",
  2637 => x"982a0772",
  2638 => x"882b87fc",
  2639 => x"80800673",
  2640 => x"982b81f0",
  2641 => x"0a067173",
  2642 => x"070780e1",
  2643 => x"800c5651",
  2644 => x"5351028c",
  2645 => x"050d0402",
  2646 => x"f8050d02",
  2647 => x"8e0580f5",
  2648 => x"2d74882b",
  2649 => x"077083ff",
  2650 => x"ff0680e1",
  2651 => x"800c5102",
  2652 => x"88050d04",
  2653 => x"02f4050d",
  2654 => x"74767853",
  2655 => x"54528071",
  2656 => x"25973872",
  2657 => x"70810554",
  2658 => x"80f52d72",
  2659 => x"70810554",
  2660 => x"81b72dff",
  2661 => x"115170eb",
  2662 => x"38807281",
  2663 => x"b72d028c",
  2664 => x"050d0402",
  2665 => x"e8050d77",
  2666 => x"56807056",
  2667 => x"54737624",
  2668 => x"b73880e9",
  2669 => x"cc08742e",
  2670 => x"af387351",
  2671 => x"80cce92d",
  2672 => x"80e18008",
  2673 => x"80e18008",
  2674 => x"09810570",
  2675 => x"80e18008",
  2676 => x"079f2a77",
  2677 => x"05811757",
  2678 => x"57535374",
  2679 => x"76248938",
  2680 => x"80e9cc08",
  2681 => x"7426d338",
  2682 => x"7280e180",
  2683 => x"0c029805",
  2684 => x"0d0402f0",
  2685 => x"050d80e0",
  2686 => x"fc081651",
  2687 => x"80d3a32d",
  2688 => x"80e18008",
  2689 => x"802ea038",
  2690 => x"8b5380e1",
  2691 => x"80085280",
  2692 => x"e7bc5180",
  2693 => x"d2f42d80",
  2694 => x"e9f80854",
  2695 => x"73802e87",
  2696 => x"3880e7bc",
  2697 => x"51732d02",
  2698 => x"90050d04",
  2699 => x"02dc050d",
  2700 => x"80705a55",
  2701 => x"7480e0fc",
  2702 => x"0825b538",
  2703 => x"80e9cc08",
  2704 => x"752ead38",
  2705 => x"785180cc",
  2706 => x"e92d80e1",
  2707 => x"80080981",
  2708 => x"057080e1",
  2709 => x"8008079f",
  2710 => x"2a760581",
  2711 => x"1b5b5654",
  2712 => x"7480e0fc",
  2713 => x"08258938",
  2714 => x"80e9cc08",
  2715 => x"7926d538",
  2716 => x"80557880",
  2717 => x"e9cc0827",
  2718 => x"81e43878",
  2719 => x"5180cce9",
  2720 => x"2d80e180",
  2721 => x"08802e81",
  2722 => x"b43880e1",
  2723 => x"80088b05",
  2724 => x"80f52d70",
  2725 => x"842a7081",
  2726 => x"06771078",
  2727 => x"842b80e7",
  2728 => x"bc0b80f5",
  2729 => x"2d5c5c53",
  2730 => x"51555673",
  2731 => x"802e80ce",
  2732 => x"38741682",
  2733 => x"2b80d782",
  2734 => x"0b80dfd0",
  2735 => x"120c5477",
  2736 => x"75311080",
  2737 => x"e9fc1155",
  2738 => x"56907470",
  2739 => x"81055681",
  2740 => x"b72da074",
  2741 => x"81b72d76",
  2742 => x"81ff0681",
  2743 => x"16585473",
  2744 => x"802e8b38",
  2745 => x"9c5380e7",
  2746 => x"bc5280d5",
  2747 => x"f5048b53",
  2748 => x"80e18008",
  2749 => x"5280e9fe",
  2750 => x"165180d6",
  2751 => x"b3047416",
  2752 => x"822b80d3",
  2753 => x"f20b80df",
  2754 => x"d0120c54",
  2755 => x"7681ff06",
  2756 => x"81165854",
  2757 => x"73802e8b",
  2758 => x"389c5380",
  2759 => x"e7bc5280",
  2760 => x"d6aa048b",
  2761 => x"5380e180",
  2762 => x"08527775",
  2763 => x"311080e9",
  2764 => x"fc055176",
  2765 => x"5580d2f4",
  2766 => x"2d80d6d2",
  2767 => x"04749029",
  2768 => x"75317010",
  2769 => x"80e9fc05",
  2770 => x"515480e1",
  2771 => x"80087481",
  2772 => x"b72d8119",
  2773 => x"59748b24",
  2774 => x"a43880d4",
  2775 => x"f2047490",
  2776 => x"29753170",
  2777 => x"1080e9fc",
  2778 => x"058c7731",
  2779 => x"57515480",
  2780 => x"7481b72d",
  2781 => x"9e14ff16",
  2782 => x"565474f3",
  2783 => x"3802a405",
  2784 => x"0d0402fc",
  2785 => x"050d80e0",
  2786 => x"fc081351",
  2787 => x"80d3a32d",
  2788 => x"80e18008",
  2789 => x"802e8a38",
  2790 => x"80e18008",
  2791 => x"5180c49d",
  2792 => x"2d800b80",
  2793 => x"e0fc0c80",
  2794 => x"d4ac2db2",
  2795 => x"9d2d0284",
  2796 => x"050d0402",
  2797 => x"fc050d72",
  2798 => x"5170fd2e",
  2799 => x"b23870fd",
  2800 => x"248b3870",
  2801 => x"fc2e80d0",
  2802 => x"3880d8a2",
  2803 => x"0470fe2e",
  2804 => x"b93870ff",
  2805 => x"2e098106",
  2806 => x"80c83880",
  2807 => x"e0fc0851",
  2808 => x"70802ebe",
  2809 => x"38ff1180",
  2810 => x"e0fc0c80",
  2811 => x"d8a20480",
  2812 => x"e0fc08f0",
  2813 => x"057080e0",
  2814 => x"fc0c5170",
  2815 => x"8025a338",
  2816 => x"800b80e0",
  2817 => x"fc0c80d8",
  2818 => x"a20480e0",
  2819 => x"fc088105",
  2820 => x"80e0fc0c",
  2821 => x"80d8a204",
  2822 => x"80e0fc08",
  2823 => x"900580e0",
  2824 => x"fc0c80d4",
  2825 => x"ac2db29d",
  2826 => x"2d028405",
  2827 => x"0d0402fc",
  2828 => x"050d800b",
  2829 => x"80e0fc0c",
  2830 => x"80d4ac2d",
  2831 => x"b1992d80",
  2832 => x"e1800880",
  2833 => x"e0ec0c80",
  2834 => x"dfc851b3",
  2835 => x"c32d0284",
  2836 => x"050d0471",
  2837 => x"80e9f80c",
  2838 => x"04000000",
  2839 => x"00ffffff",
  2840 => x"ff00ffff",
  2841 => x"ffff00ff",
  2842 => x"ffffff00",
  2843 => x"30313233",
  2844 => x"34353637",
  2845 => x"38394142",
  2846 => x"43444546",
  2847 => x"00000000",
  2848 => x"52657365",
  2849 => x"74000000",
  2850 => x"5363616e",
  2851 => x"6c696e65",
  2852 => x"73000000",
  2853 => x"50414c20",
  2854 => x"2f204e54",
  2855 => x"53430000",
  2856 => x"436f6c6f",
  2857 => x"72000000",
  2858 => x"44696666",
  2859 => x"6963756c",
  2860 => x"74792041",
  2861 => x"00000000",
  2862 => x"44696666",
  2863 => x"6963756c",
  2864 => x"74792042",
  2865 => x"00000000",
  2866 => x"2a537570",
  2867 => x"65726368",
  2868 => x"69702069",
  2869 => x"6e206361",
  2870 => x"72747269",
  2871 => x"64676500",
  2872 => x"2a42616e",
  2873 => x"6b204530",
  2874 => x"00000000",
  2875 => x"2a42616e",
  2876 => x"6b204537",
  2877 => x"00000000",
  2878 => x"53656c65",
  2879 => x"63740000",
  2880 => x"53746172",
  2881 => x"74000000",
  2882 => x"4c6f6164",
  2883 => x"20524f4d",
  2884 => x"20100000",
  2885 => x"45786974",
  2886 => x"00000000",
  2887 => x"524f4d20",
  2888 => x"6c6f6164",
  2889 => x"696e6720",
  2890 => x"6661696c",
  2891 => x"65640000",
  2892 => x"4f4b0000",
  2893 => x"496e6974",
  2894 => x"69616c69",
  2895 => x"7a696e67",
  2896 => x"20534420",
  2897 => x"63617264",
  2898 => x"0a000000",
  2899 => x"436f6c6c",
  2900 => x"6563746f",
  2901 => x"72566973",
  2902 => x"696f6e00",
  2903 => x"64626732",
  2904 => x"00000000",
  2905 => x"16200000",
  2906 => x"14200000",
  2907 => x"15200000",
  2908 => x"53442069",
  2909 => x"6e69742e",
  2910 => x"2e2e0a00",
  2911 => x"53442063",
  2912 => x"61726420",
  2913 => x"72657365",
  2914 => x"74206661",
  2915 => x"696c6564",
  2916 => x"210a0000",
  2917 => x"53444843",
  2918 => x"20657272",
  2919 => x"6f72210a",
  2920 => x"00000000",
  2921 => x"57726974",
  2922 => x"65206661",
  2923 => x"696c6564",
  2924 => x"0a000000",
  2925 => x"52656164",
  2926 => x"20666169",
  2927 => x"6c65640a",
  2928 => x"00000000",
  2929 => x"43617264",
  2930 => x"20696e69",
  2931 => x"74206661",
  2932 => x"696c6564",
  2933 => x"0a000000",
  2934 => x"46415431",
  2935 => x"36202020",
  2936 => x"00000000",
  2937 => x"46415433",
  2938 => x"32202020",
  2939 => x"00000000",
  2940 => x"4e6f2070",
  2941 => x"61727469",
  2942 => x"74696f6e",
  2943 => x"20736967",
  2944 => x"0a000000",
  2945 => x"42616420",
  2946 => x"70617274",
  2947 => x"0a000000",
  2948 => x"4261636b",
  2949 => x"00000000",
  2950 => x"00000002",
  2951 => x"00002c6c",
  2952 => x"00003130",
  2953 => x"00000002",
  2954 => x"000030a8",
  2955 => x"0000140a",
  2956 => x"00000002",
  2957 => x"000030ec",
  2958 => x"00001326",
  2959 => x"00000002",
  2960 => x"00002c80",
  2961 => x"0000035a",
  2962 => x"00000001",
  2963 => x"00002c88",
  2964 => x"00000000",
  2965 => x"00000001",
  2966 => x"00002c94",
  2967 => x"00000001",
  2968 => x"00000001",
  2969 => x"00002ca0",
  2970 => x"00000002",
  2971 => x"00000001",
  2972 => x"00002ca8",
  2973 => x"00000003",
  2974 => x"00000001",
  2975 => x"00002cb8",
  2976 => x"00000004",
  2977 => x"00000001",
  2978 => x"00002cc8",
  2979 => x"00000005",
  2980 => x"00000001",
  2981 => x"00002ce0",
  2982 => x"00000008",
  2983 => x"00000001",
  2984 => x"00002cec",
  2985 => x"00000009",
  2986 => x"00000002",
  2987 => x"00002cf8",
  2988 => x"0000036e",
  2989 => x"00000002",
  2990 => x"00002d00",
  2991 => x"00000a3f",
  2992 => x"00000002",
  2993 => x"00002d08",
  2994 => x"00002c2e",
  2995 => x"00000002",
  2996 => x"00002d14",
  2997 => x"000018b6",
  2998 => x"00000000",
  2999 => x"00000000",
  3000 => x"00000000",
  3001 => x"00000004",
  3002 => x"00002d1c",
  3003 => x"00002ee4",
  3004 => x"00000004",
  3005 => x"00002d30",
  3006 => x"00002e24",
  3007 => x"00000000",
  3008 => x"00000000",
  3009 => x"00000000",
  3010 => x"00000000",
  3011 => x"00000000",
  3012 => x"00000000",
  3013 => x"00000000",
  3014 => x"00000000",
  3015 => x"00000000",
  3016 => x"00000000",
  3017 => x"00000000",
  3018 => x"00000000",
  3019 => x"00000000",
  3020 => x"00000000",
  3021 => x"00000000",
  3022 => x"00000000",
  3023 => x"00000000",
  3024 => x"00000000",
  3025 => x"00000000",
  3026 => x"00000000",
  3027 => x"761c1c1c",
  3028 => x"1c1c051c",
  3029 => x"1c1c1c1c",
  3030 => x"f2f5ebf4",
  3031 => x"5a000000",
  3032 => x"00000000",
  3033 => x"00000000",
  3034 => x"00000000",
  3035 => x"00000000",
  3036 => x"00000000",
  3037 => x"00000000",
  3038 => x"00000000",
  3039 => x"00000000",
  3040 => x"00000000",
  3041 => x"00000000",
  3042 => x"00000000",
  3043 => x"00000000",
  3044 => x"00000000",
  3045 => x"00000000",
  3046 => x"00000000",
  3047 => x"00000000",
  3048 => x"00000000",
  3049 => x"00000000",
  3050 => x"0001ffff",
  3051 => x"0001ffff",
  3052 => x"0001ffff",
  3053 => x"00000000",
  3054 => x"00000000",
  3055 => x"00000006",
  3056 => x"00000000",
  3057 => x"00000000",
  3058 => x"00000002",
  3059 => x"000034fc",
  3060 => x"000029f2",
  3061 => x"00000002",
  3062 => x"0000351a",
  3063 => x"000029f2",
  3064 => x"00000002",
  3065 => x"00003538",
  3066 => x"000029f2",
  3067 => x"00000002",
  3068 => x"00003556",
  3069 => x"000029f2",
  3070 => x"00000002",
  3071 => x"00003574",
  3072 => x"000029f2",
  3073 => x"00000002",
  3074 => x"00003592",
  3075 => x"000029f2",
  3076 => x"00000002",
  3077 => x"000035b0",
  3078 => x"000029f2",
  3079 => x"00000002",
  3080 => x"000035ce",
  3081 => x"000029f2",
  3082 => x"00000002",
  3083 => x"000035ec",
  3084 => x"000029f2",
  3085 => x"00000002",
  3086 => x"0000360a",
  3087 => x"000029f2",
  3088 => x"00000002",
  3089 => x"00003628",
  3090 => x"000029f2",
  3091 => x"00000002",
  3092 => x"00003646",
  3093 => x"000029f2",
  3094 => x"00000002",
  3095 => x"00003664",
  3096 => x"000029f2",
  3097 => x"00000004",
  3098 => x"00002e10",
  3099 => x"00000000",
  3100 => x"00000000",
  3101 => x"00000000",
  3102 => x"00002bb3",
  3103 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

