-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80dd",
     9 => x"a0080b0b",
    10 => x"80dda408",
    11 => x"0b0b80dd",
    12 => x"a8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"dda80c0b",
    16 => x"0b80dda4",
    17 => x"0c0b0b80",
    18 => x"dda00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d5b8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80dda070",
    57 => x"80e7d827",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a6b7",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80dd",
    65 => x"b00c9f0b",
    66 => x"80ddb40c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"ddb408ff",
    70 => x"0580ddb4",
    71 => x"0c80ddb4",
    72 => x"088025e8",
    73 => x"3880ddb0",
    74 => x"08ff0580",
    75 => x"ddb00c80",
    76 => x"ddb00880",
    77 => x"25d03880",
    78 => x"0b80ddb4",
    79 => x"0c800b80",
    80 => x"ddb00c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80ddb008",
   100 => x"25913882",
   101 => x"c82d80dd",
   102 => x"b008ff05",
   103 => x"80ddb00c",
   104 => x"838a0480",
   105 => x"ddb00880",
   106 => x"ddb40853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80ddb008",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"ddb40881",
   116 => x"0580ddb4",
   117 => x"0c80ddb4",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80ddb4",
   121 => x"0c80ddb0",
   122 => x"08810580",
   123 => x"ddb00c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480dd",
   128 => x"b4088105",
   129 => x"80ddb40c",
   130 => x"80ddb408",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80ddb4",
   134 => x"0c80ddb0",
   135 => x"08810580",
   136 => x"ddb00c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"ddb80cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"ddb80c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280dd",
   177 => x"b8088407",
   178 => x"80ddb80c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80d8",
   183 => x"dc0c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80ddb8",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80dd",
   208 => x"a00c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02f4050d",
  1093 => x"80d8f40b",
  1094 => x"80f52d80",
  1095 => x"dbdc0870",
  1096 => x"81065354",
  1097 => x"5270802e",
  1098 => x"85387184",
  1099 => x"07527281",
  1100 => x"2a708106",
  1101 => x"51517080",
  1102 => x"2e853871",
  1103 => x"82075272",
  1104 => x"822a7081",
  1105 => x"06515170",
  1106 => x"802e8538",
  1107 => x"71810752",
  1108 => x"72832a70",
  1109 => x"81065151",
  1110 => x"70802e85",
  1111 => x"38718807",
  1112 => x"5272842a",
  1113 => x"70810651",
  1114 => x"5170802e",
  1115 => x"85387190",
  1116 => x"07527285",
  1117 => x"2a708106",
  1118 => x"51517080",
  1119 => x"2e853871",
  1120 => x"a0075272",
  1121 => x"882a7081",
  1122 => x"06515170",
  1123 => x"802e8638",
  1124 => x"7180c007",
  1125 => x"5272892a",
  1126 => x"70810651",
  1127 => x"5170802e",
  1128 => x"86387181",
  1129 => x"80075271",
  1130 => x"fc0c7180",
  1131 => x"dda00c02",
  1132 => x"8c050d04",
  1133 => x"02cc050d",
  1134 => x"7e5d800b",
  1135 => x"80dbdc08",
  1136 => x"81800671",
  1137 => x"5c5d5b81",
  1138 => x"0bec0c84",
  1139 => x"0bec0c7c",
  1140 => x"5280ddbc",
  1141 => x"5180cc87",
  1142 => x"2d80dda0",
  1143 => x"087b2e80",
  1144 => x"ff3880dd",
  1145 => x"c0087bff",
  1146 => x"12575957",
  1147 => x"747b2e8b",
  1148 => x"38811875",
  1149 => x"812a5658",
  1150 => x"74f738f7",
  1151 => x"1858815b",
  1152 => x"80772580",
  1153 => x"db387752",
  1154 => x"745184a8",
  1155 => x"2d80de90",
  1156 => x"5280ddbc",
  1157 => x"5180cedc",
  1158 => x"2d80dda0",
  1159 => x"08802ea6",
  1160 => x"3880de90",
  1161 => x"597ba738",
  1162 => x"83ff5678",
  1163 => x"7081055a",
  1164 => x"80f52d7a",
  1165 => x"811c5ce4",
  1166 => x"0ce80cff",
  1167 => x"16567580",
  1168 => x"25e938a4",
  1169 => x"ce0480dd",
  1170 => x"a0085b84",
  1171 => x"805780dd",
  1172 => x"bc5180ce",
  1173 => x"ab2dfc80",
  1174 => x"17811656",
  1175 => x"57a48004",
  1176 => x"80ddc008",
  1177 => x"f80c881d",
  1178 => x"55807580",
  1179 => x"f52d7081",
  1180 => x"ff065558",
  1181 => x"5472742e",
  1182 => x"b6388115",
  1183 => x"80f52d53",
  1184 => x"72742eab",
  1185 => x"38738216",
  1186 => x"80f52d54",
  1187 => x"567280d3",
  1188 => x"2e098106",
  1189 => x"83388156",
  1190 => x"7280f332",
  1191 => x"70098105",
  1192 => x"70802578",
  1193 => x"07515153",
  1194 => x"72802e83",
  1195 => x"38a05480",
  1196 => x"7781ff06",
  1197 => x"54567280",
  1198 => x"c52e0981",
  1199 => x"06833881",
  1200 => x"567280e5",
  1201 => x"32700981",
  1202 => x"05708025",
  1203 => x"78075151",
  1204 => x"5372802e",
  1205 => x"a4388115",
  1206 => x"80f52d53",
  1207 => x"72b02e09",
  1208 => x"81068938",
  1209 => x"73828007",
  1210 => x"54a5f904",
  1211 => x"72b72e09",
  1212 => x"81068638",
  1213 => x"73848007",
  1214 => x"5473802e",
  1215 => x"913880db",
  1216 => x"dc08f9df",
  1217 => x"06740780",
  1218 => x"dbdc0ca2",
  1219 => x"902d810b",
  1220 => x"e00c8051",
  1221 => x"86da2d86",
  1222 => x"c72d7a80",
  1223 => x"2e883880",
  1224 => x"d8e051a6",
  1225 => x"aa0480da",
  1226 => x"8851b0ae",
  1227 => x"2d7a80dd",
  1228 => x"a00c02b4",
  1229 => x"050d0402",
  1230 => x"f4050d84",
  1231 => x"0bec0cad",
  1232 => x"eb2da7c5",
  1233 => x"2d81f92d",
  1234 => x"8352adce",
  1235 => x"2d815185",
  1236 => x"8d2dff12",
  1237 => x"52718025",
  1238 => x"f138840b",
  1239 => x"ec0c80d7",
  1240 => x"905186a0",
  1241 => x"2d80c2ac",
  1242 => x"2d80dda0",
  1243 => x"08802ebe",
  1244 => x"38a3b451",
  1245 => x"80d5b22d",
  1246 => x"80d8e051",
  1247 => x"b0ae2dae",
  1248 => x"8d2da8f0",
  1249 => x"2d80dda0",
  1250 => x"08810652",
  1251 => x"71802e86",
  1252 => x"38805194",
  1253 => x"bf2db0c1",
  1254 => x"2d80dda0",
  1255 => x"0852a290",
  1256 => x"2d865371",
  1257 => x"83388453",
  1258 => x"72ec0ca7",
  1259 => x"8204800b",
  1260 => x"80dda00c",
  1261 => x"028c050d",
  1262 => x"0471980c",
  1263 => x"04ffb008",
  1264 => x"80dda00c",
  1265 => x"04810bff",
  1266 => x"b00c0480",
  1267 => x"0bffb00c",
  1268 => x"0402d805",
  1269 => x"0dffb408",
  1270 => x"87ffff06",
  1271 => x"5a815480",
  1272 => x"7080dbc8",
  1273 => x"0880dbcc",
  1274 => x"0880dba4",
  1275 => x"5b59575a",
  1276 => x"58797406",
  1277 => x"75750652",
  1278 => x"5271712e",
  1279 => x"8d388077",
  1280 => x"818a2d73",
  1281 => x"09750672",
  1282 => x"07557680",
  1283 => x"e02d7083",
  1284 => x"ffff0653",
  1285 => x"517180e4",
  1286 => x"2e098106",
  1287 => x"a2387474",
  1288 => x"06707776",
  1289 => x"06327009",
  1290 => x"81057072",
  1291 => x"079f2a7b",
  1292 => x"0577097a",
  1293 => x"0674075a",
  1294 => x"5b535353",
  1295 => x"a8cd0471",
  1296 => x"80e42689",
  1297 => x"38811151",
  1298 => x"7077818a",
  1299 => x"2d731081",
  1300 => x"1a821959",
  1301 => x"5a549079",
  1302 => x"25ff9638",
  1303 => x"7580dbcc",
  1304 => x"0c7480db",
  1305 => x"c80c7780",
  1306 => x"dda00c02",
  1307 => x"a8050d04",
  1308 => x"02d0050d",
  1309 => x"805caa80",
  1310 => x"0480dda0",
  1311 => x"0881f02e",
  1312 => x"0981068a",
  1313 => x"38810b80",
  1314 => x"dbd40caa",
  1315 => x"800480dd",
  1316 => x"a00881e0",
  1317 => x"2e098106",
  1318 => x"8a38810b",
  1319 => x"80dbd80c",
  1320 => x"aa800480",
  1321 => x"dda00852",
  1322 => x"80dbd808",
  1323 => x"802e8938",
  1324 => x"80dda008",
  1325 => x"81800552",
  1326 => x"71842c72",
  1327 => x"8f065353",
  1328 => x"80dbd408",
  1329 => x"802e9a38",
  1330 => x"72842980",
  1331 => x"daac0572",
  1332 => x"1381712b",
  1333 => x"70097308",
  1334 => x"06730c51",
  1335 => x"5353a9f4",
  1336 => x"04728429",
  1337 => x"80daac05",
  1338 => x"72138371",
  1339 => x"2b720807",
  1340 => x"720c5353",
  1341 => x"800b80db",
  1342 => x"d80c800b",
  1343 => x"80dbd40c",
  1344 => x"80ddc851",
  1345 => x"acc12d80",
  1346 => x"dda008ff",
  1347 => x"24feea38",
  1348 => x"a7d12d80",
  1349 => x"dda00880",
  1350 => x"2e81b038",
  1351 => x"8159800b",
  1352 => x"80dbd008",
  1353 => x"80dbcc08",
  1354 => x"80db805a",
  1355 => x"5c5c587a",
  1356 => x"79067a7a",
  1357 => x"06545271",
  1358 => x"732e80f8",
  1359 => x"38720981",
  1360 => x"05707407",
  1361 => x"802580da",
  1362 => x"ec1a80f5",
  1363 => x"2d70842c",
  1364 => x"718f0658",
  1365 => x"53575752",
  1366 => x"75802ea3",
  1367 => x"38718429",
  1368 => x"80daac05",
  1369 => x"74158371",
  1370 => x"2b720807",
  1371 => x"720c5452",
  1372 => x"7680e02d",
  1373 => x"81055271",
  1374 => x"77818a2d",
  1375 => x"ab950471",
  1376 => x"842980da",
  1377 => x"ac057415",
  1378 => x"81712b70",
  1379 => x"09730806",
  1380 => x"730c5153",
  1381 => x"53748532",
  1382 => x"70098105",
  1383 => x"70802551",
  1384 => x"51527580",
  1385 => x"2e8e3881",
  1386 => x"70730653",
  1387 => x"5371802e",
  1388 => x"8338725c",
  1389 => x"78108119",
  1390 => x"82195959",
  1391 => x"59907825",
  1392 => x"feed3880",
  1393 => x"dbcc0880",
  1394 => x"dbd00c7b",
  1395 => x"80dda00c",
  1396 => x"02b0050d",
  1397 => x"0402f805",
  1398 => x"0d80daac",
  1399 => x"528f5180",
  1400 => x"72708405",
  1401 => x"540cff11",
  1402 => x"51708025",
  1403 => x"f2380288",
  1404 => x"050d0402",
  1405 => x"f0050d75",
  1406 => x"51a7cb2d",
  1407 => x"70822cfc",
  1408 => x"0680daac",
  1409 => x"1172109e",
  1410 => x"06710870",
  1411 => x"722a7083",
  1412 => x"0682742b",
  1413 => x"70097406",
  1414 => x"760c5451",
  1415 => x"56575351",
  1416 => x"53a7c52d",
  1417 => x"7180dda0",
  1418 => x"0c029005",
  1419 => x"0d0402fc",
  1420 => x"050d7251",
  1421 => x"80710c80",
  1422 => x"0b84120c",
  1423 => x"0284050d",
  1424 => x"0402f005",
  1425 => x"0d757008",
  1426 => x"84120853",
  1427 => x"5353ff54",
  1428 => x"71712ea8",
  1429 => x"38a7cb2d",
  1430 => x"84130870",
  1431 => x"84291488",
  1432 => x"11700870",
  1433 => x"81ff0684",
  1434 => x"18088111",
  1435 => x"8706841a",
  1436 => x"0c535155",
  1437 => x"515151a7",
  1438 => x"c52d7154",
  1439 => x"7380dda0",
  1440 => x"0c029005",
  1441 => x"0d0402f8",
  1442 => x"050da7cb",
  1443 => x"2de00870",
  1444 => x"8b2a7081",
  1445 => x"06515252",
  1446 => x"70802ea1",
  1447 => x"3880ddc8",
  1448 => x"08708429",
  1449 => x"80ddd005",
  1450 => x"7381ff06",
  1451 => x"710c5151",
  1452 => x"80ddc808",
  1453 => x"81118706",
  1454 => x"80ddc80c",
  1455 => x"51800b80",
  1456 => x"ddf00ca7",
  1457 => x"bd2da7c5",
  1458 => x"2d028805",
  1459 => x"0d0402fc",
  1460 => x"050da7cb",
  1461 => x"2d810b80",
  1462 => x"ddf00ca7",
  1463 => x"c52d80dd",
  1464 => x"f0085170",
  1465 => x"f9380284",
  1466 => x"050d0402",
  1467 => x"fc050d80",
  1468 => x"ddc851ac",
  1469 => x"ae2dabd5",
  1470 => x"2dad8651",
  1471 => x"a7b92d02",
  1472 => x"84050d04",
  1473 => x"80ddfc08",
  1474 => x"80dda00c",
  1475 => x"0402fc05",
  1476 => x"0d810b80",
  1477 => x"dbe00c81",
  1478 => x"51858d2d",
  1479 => x"0284050d",
  1480 => x"0402fc05",
  1481 => x"0daeab04",
  1482 => x"a8f02d80",
  1483 => x"f651abf3",
  1484 => x"2d80dda0",
  1485 => x"08f23880",
  1486 => x"da51abf3",
  1487 => x"2d80dda0",
  1488 => x"08e63880",
  1489 => x"dda00880",
  1490 => x"dbe00c80",
  1491 => x"dda00851",
  1492 => x"858d2d02",
  1493 => x"84050d04",
  1494 => x"02ec050d",
  1495 => x"76548052",
  1496 => x"870b8815",
  1497 => x"80f52d56",
  1498 => x"53747224",
  1499 => x"8338a053",
  1500 => x"72518384",
  1501 => x"2d81128b",
  1502 => x"1580f52d",
  1503 => x"54527272",
  1504 => x"25de3802",
  1505 => x"94050d04",
  1506 => x"02f0050d",
  1507 => x"80ddfc08",
  1508 => x"5481f92d",
  1509 => x"800b80de",
  1510 => x"800c7308",
  1511 => x"802e8189",
  1512 => x"38820b80",
  1513 => x"ddb40c80",
  1514 => x"de80088f",
  1515 => x"0680ddb0",
  1516 => x"0c730852",
  1517 => x"71832e96",
  1518 => x"38718326",
  1519 => x"89387181",
  1520 => x"2eb038b0",
  1521 => x"92047185",
  1522 => x"2ea038b0",
  1523 => x"92048814",
  1524 => x"80f52d84",
  1525 => x"150880d7",
  1526 => x"a8535452",
  1527 => x"86a02d71",
  1528 => x"84291370",
  1529 => x"085252b0",
  1530 => x"96047351",
  1531 => x"aed82db0",
  1532 => x"920480db",
  1533 => x"dc088815",
  1534 => x"082c7081",
  1535 => x"06515271",
  1536 => x"802e8838",
  1537 => x"80d7ac51",
  1538 => x"b08f0480",
  1539 => x"d7b05186",
  1540 => x"a02d8414",
  1541 => x"085186a0",
  1542 => x"2d80de80",
  1543 => x"08810580",
  1544 => x"de800c8c",
  1545 => x"1454af9a",
  1546 => x"04029005",
  1547 => x"0d047180",
  1548 => x"ddfc0caf",
  1549 => x"882d80de",
  1550 => x"8008ff05",
  1551 => x"80de840c",
  1552 => x"0402e805",
  1553 => x"0d80ddfc",
  1554 => x"0880de88",
  1555 => x"08575580",
  1556 => x"f651abf3",
  1557 => x"2d80dda0",
  1558 => x"08812a70",
  1559 => x"81065152",
  1560 => x"71802ea4",
  1561 => x"38b0eb04",
  1562 => x"a8f02d80",
  1563 => x"f651abf3",
  1564 => x"2d80dda0",
  1565 => x"08f23880",
  1566 => x"dbe00881",
  1567 => x"327080db",
  1568 => x"e00c7052",
  1569 => x"52858d2d",
  1570 => x"800b80dd",
  1571 => x"f40c800b",
  1572 => x"80ddf80c",
  1573 => x"80dbe008",
  1574 => x"838d3880",
  1575 => x"da51abf3",
  1576 => x"2d80dda0",
  1577 => x"08802e8c",
  1578 => x"3880ddf4",
  1579 => x"08818007",
  1580 => x"80ddf40c",
  1581 => x"80d951ab",
  1582 => x"f32d80dd",
  1583 => x"a008802e",
  1584 => x"8c3880dd",
  1585 => x"f40880c0",
  1586 => x"0780ddf4",
  1587 => x"0c819451",
  1588 => x"abf32d80",
  1589 => x"dda00880",
  1590 => x"2e8b3880",
  1591 => x"ddf40890",
  1592 => x"0780ddf4",
  1593 => x"0c819151",
  1594 => x"abf32d80",
  1595 => x"dda00880",
  1596 => x"2e8b3880",
  1597 => x"ddf408a0",
  1598 => x"0780ddf4",
  1599 => x"0c81f551",
  1600 => x"abf32d80",
  1601 => x"dda00880",
  1602 => x"2e8b3880",
  1603 => x"ddf40881",
  1604 => x"0780ddf4",
  1605 => x"0c81f251",
  1606 => x"abf32d80",
  1607 => x"dda00880",
  1608 => x"2e8b3880",
  1609 => x"ddf40882",
  1610 => x"0780ddf4",
  1611 => x"0c81eb51",
  1612 => x"abf32d80",
  1613 => x"dda00880",
  1614 => x"2e8b3880",
  1615 => x"ddf40884",
  1616 => x"0780ddf4",
  1617 => x"0c81f451",
  1618 => x"abf32d80",
  1619 => x"dda00880",
  1620 => x"2e8b3880",
  1621 => x"ddf40888",
  1622 => x"0780ddf4",
  1623 => x"0c80d851",
  1624 => x"abf32d80",
  1625 => x"dda00880",
  1626 => x"2e8c3880",
  1627 => x"ddf80881",
  1628 => x"800780dd",
  1629 => x"f80c9251",
  1630 => x"abf32d80",
  1631 => x"dda00880",
  1632 => x"2e8c3880",
  1633 => x"ddf80880",
  1634 => x"c00780dd",
  1635 => x"f80c9451",
  1636 => x"abf32d80",
  1637 => x"dda00880",
  1638 => x"2e8b3880",
  1639 => x"ddf80890",
  1640 => x"0780ddf8",
  1641 => x"0c9151ab",
  1642 => x"f32d80dd",
  1643 => x"a008802e",
  1644 => x"8b3880dd",
  1645 => x"f808a007",
  1646 => x"80ddf80c",
  1647 => x"9d51abf3",
  1648 => x"2d80dda0",
  1649 => x"08802e8b",
  1650 => x"3880ddf8",
  1651 => x"08810780",
  1652 => x"ddf80c9b",
  1653 => x"51abf32d",
  1654 => x"80dda008",
  1655 => x"802e8b38",
  1656 => x"80ddf808",
  1657 => x"820780dd",
  1658 => x"f80c9c51",
  1659 => x"abf32d80",
  1660 => x"dda00880",
  1661 => x"2e8b3880",
  1662 => x"ddf80884",
  1663 => x"0780ddf8",
  1664 => x"0ca351ab",
  1665 => x"f32d80dd",
  1666 => x"a008802e",
  1667 => x"8b3880dd",
  1668 => x"f8088807",
  1669 => x"80ddf80c",
  1670 => x"81fd51ab",
  1671 => x"f32d81fa",
  1672 => x"51abf32d",
  1673 => x"b9fc0481",
  1674 => x"f551abf3",
  1675 => x"2d80dda0",
  1676 => x"08812a70",
  1677 => x"81065152",
  1678 => x"71802eb3",
  1679 => x"3880de84",
  1680 => x"08527180",
  1681 => x"2e8a38ff",
  1682 => x"1280de84",
  1683 => x"0cb4ef04",
  1684 => x"80de8008",
  1685 => x"1080de80",
  1686 => x"08057084",
  1687 => x"29165152",
  1688 => x"88120880",
  1689 => x"2e8938ff",
  1690 => x"51881208",
  1691 => x"52712d81",
  1692 => x"f251abf3",
  1693 => x"2d80dda0",
  1694 => x"08812a70",
  1695 => x"81065152",
  1696 => x"71802eb4",
  1697 => x"3880de80",
  1698 => x"08ff1180",
  1699 => x"de840856",
  1700 => x"53537372",
  1701 => x"258a3881",
  1702 => x"1480de84",
  1703 => x"0cb5b804",
  1704 => x"72101370",
  1705 => x"84291651",
  1706 => x"52881208",
  1707 => x"802e8938",
  1708 => x"fe518812",
  1709 => x"0852712d",
  1710 => x"81fd51ab",
  1711 => x"f32d80dd",
  1712 => x"a008812a",
  1713 => x"70810651",
  1714 => x"5271802e",
  1715 => x"b13880de",
  1716 => x"8408802e",
  1717 => x"8a38800b",
  1718 => x"80de840c",
  1719 => x"b5fe0480",
  1720 => x"de800810",
  1721 => x"80de8008",
  1722 => x"05708429",
  1723 => x"16515288",
  1724 => x"1208802e",
  1725 => x"8938fd51",
  1726 => x"88120852",
  1727 => x"712d81fa",
  1728 => x"51abf32d",
  1729 => x"80dda008",
  1730 => x"812a7081",
  1731 => x"06515271",
  1732 => x"802eb138",
  1733 => x"80de8008",
  1734 => x"ff115452",
  1735 => x"80de8408",
  1736 => x"73258938",
  1737 => x"7280de84",
  1738 => x"0cb6c404",
  1739 => x"71101270",
  1740 => x"84291651",
  1741 => x"52881208",
  1742 => x"802e8938",
  1743 => x"fc518812",
  1744 => x"0852712d",
  1745 => x"80de8408",
  1746 => x"70535473",
  1747 => x"802e8a38",
  1748 => x"8c15ff15",
  1749 => x"5555b6cb",
  1750 => x"04820b80",
  1751 => x"ddb40c71",
  1752 => x"8f0680dd",
  1753 => x"b00c81eb",
  1754 => x"51abf32d",
  1755 => x"80dda008",
  1756 => x"812a7081",
  1757 => x"06515271",
  1758 => x"802ead38",
  1759 => x"7408852e",
  1760 => x"098106a4",
  1761 => x"38881580",
  1762 => x"f52dff05",
  1763 => x"52718816",
  1764 => x"81b72d71",
  1765 => x"982b5271",
  1766 => x"80258838",
  1767 => x"800b8816",
  1768 => x"81b72d74",
  1769 => x"51aed82d",
  1770 => x"81f451ab",
  1771 => x"f32d80dd",
  1772 => x"a008812a",
  1773 => x"70810651",
  1774 => x"5271802e",
  1775 => x"b3387408",
  1776 => x"852e0981",
  1777 => x"06aa3888",
  1778 => x"1580f52d",
  1779 => x"81055271",
  1780 => x"881681b7",
  1781 => x"2d7181ff",
  1782 => x"068b1680",
  1783 => x"f52d5452",
  1784 => x"72722787",
  1785 => x"38728816",
  1786 => x"81b72d74",
  1787 => x"51aed82d",
  1788 => x"80da51ab",
  1789 => x"f32d80dd",
  1790 => x"a008812a",
  1791 => x"70810651",
  1792 => x"5271802e",
  1793 => x"81ad3880",
  1794 => x"ddfc0880",
  1795 => x"de840855",
  1796 => x"5373802e",
  1797 => x"8a388c13",
  1798 => x"ff155553",
  1799 => x"b8910472",
  1800 => x"08527182",
  1801 => x"2ea63871",
  1802 => x"82268938",
  1803 => x"71812eaa",
  1804 => x"38b9b304",
  1805 => x"71832eb4",
  1806 => x"3871842e",
  1807 => x"09810680",
  1808 => x"f2388813",
  1809 => x"0851b0ae",
  1810 => x"2db9b304",
  1811 => x"80de8408",
  1812 => x"51881308",
  1813 => x"52712db9",
  1814 => x"b304810b",
  1815 => x"8814082b",
  1816 => x"80dbdc08",
  1817 => x"3280dbdc",
  1818 => x"0cb98704",
  1819 => x"881380f5",
  1820 => x"2d81058b",
  1821 => x"1480f52d",
  1822 => x"53547174",
  1823 => x"24833880",
  1824 => x"54738814",
  1825 => x"81b72daf",
  1826 => x"882db9b3",
  1827 => x"04750880",
  1828 => x"2ea43875",
  1829 => x"0851abf3",
  1830 => x"2d80dda0",
  1831 => x"08810652",
  1832 => x"71802e8c",
  1833 => x"3880de84",
  1834 => x"08518416",
  1835 => x"0852712d",
  1836 => x"88165675",
  1837 => x"d8388054",
  1838 => x"800b80dd",
  1839 => x"b40c738f",
  1840 => x"0680ddb0",
  1841 => x"0ca05273",
  1842 => x"80de8408",
  1843 => x"2e098106",
  1844 => x"993880de",
  1845 => x"8008ff05",
  1846 => x"74327009",
  1847 => x"81057072",
  1848 => x"079f2a91",
  1849 => x"71315151",
  1850 => x"53537151",
  1851 => x"83842d81",
  1852 => x"14548e74",
  1853 => x"25c23880",
  1854 => x"dbe00852",
  1855 => x"7180dda0",
  1856 => x"0c029805",
  1857 => x"0d0402f4",
  1858 => x"050dd452",
  1859 => x"81ff720c",
  1860 => x"71085381",
  1861 => x"ff720c72",
  1862 => x"882b83fe",
  1863 => x"80067208",
  1864 => x"7081ff06",
  1865 => x"51525381",
  1866 => x"ff720c72",
  1867 => x"7107882b",
  1868 => x"72087081",
  1869 => x"ff065152",
  1870 => x"5381ff72",
  1871 => x"0c727107",
  1872 => x"882b7208",
  1873 => x"7081ff06",
  1874 => x"720780dd",
  1875 => x"a00c5253",
  1876 => x"028c050d",
  1877 => x"0402f405",
  1878 => x"0d747671",
  1879 => x"81ff06d4",
  1880 => x"0c535380",
  1881 => x"de8c0885",
  1882 => x"3871892b",
  1883 => x"5271982a",
  1884 => x"d40c7190",
  1885 => x"2a7081ff",
  1886 => x"06d40c51",
  1887 => x"71882a70",
  1888 => x"81ff06d4",
  1889 => x"0c517181",
  1890 => x"ff06d40c",
  1891 => x"72902a70",
  1892 => x"81ff06d4",
  1893 => x"0c51d408",
  1894 => x"7081ff06",
  1895 => x"515182b8",
  1896 => x"bf527081",
  1897 => x"ff2e0981",
  1898 => x"06943881",
  1899 => x"ff0bd40c",
  1900 => x"d4087081",
  1901 => x"ff06ff14",
  1902 => x"54515171",
  1903 => x"e5387080",
  1904 => x"dda00c02",
  1905 => x"8c050d04",
  1906 => x"02fc050d",
  1907 => x"81c75181",
  1908 => x"ff0bd40c",
  1909 => x"ff115170",
  1910 => x"8025f438",
  1911 => x"0284050d",
  1912 => x"0402f405",
  1913 => x"0d81ff0b",
  1914 => x"d40c9353",
  1915 => x"805287fc",
  1916 => x"80c151ba",
  1917 => x"d52d80dd",
  1918 => x"a0088b38",
  1919 => x"81ff0bd4",
  1920 => x"0c8153bc",
  1921 => x"8f04bbc8",
  1922 => x"2dff1353",
  1923 => x"72de3872",
  1924 => x"80dda00c",
  1925 => x"028c050d",
  1926 => x"0402ec05",
  1927 => x"0d810b80",
  1928 => x"de8c0c84",
  1929 => x"54d00870",
  1930 => x"8f2a7081",
  1931 => x"06515153",
  1932 => x"72f33872",
  1933 => x"d00cbbc8",
  1934 => x"2d80d7b4",
  1935 => x"5186a02d",
  1936 => x"d008708f",
  1937 => x"2a708106",
  1938 => x"51515372",
  1939 => x"f338810b",
  1940 => x"d00cb153",
  1941 => x"805284d4",
  1942 => x"80c051ba",
  1943 => x"d52d80dd",
  1944 => x"a008812e",
  1945 => x"93387282",
  1946 => x"2ebf38ff",
  1947 => x"135372e4",
  1948 => x"38ff1454",
  1949 => x"73ffae38",
  1950 => x"bbc82d83",
  1951 => x"aa52849c",
  1952 => x"80c851ba",
  1953 => x"d52d80dd",
  1954 => x"a008812e",
  1955 => x"09810693",
  1956 => x"38ba862d",
  1957 => x"80dda008",
  1958 => x"83ffff06",
  1959 => x"537283aa",
  1960 => x"2e9f38bb",
  1961 => x"e12dbdbc",
  1962 => x"0480d7c0",
  1963 => x"5186a02d",
  1964 => x"8053bf91",
  1965 => x"0480d7d8",
  1966 => x"5186a02d",
  1967 => x"8054bee2",
  1968 => x"0481ff0b",
  1969 => x"d40cb154",
  1970 => x"bbc82d8f",
  1971 => x"cf538052",
  1972 => x"87fc80f7",
  1973 => x"51bad52d",
  1974 => x"80dda008",
  1975 => x"5580dda0",
  1976 => x"08812e09",
  1977 => x"81069c38",
  1978 => x"81ff0bd4",
  1979 => x"0c820a52",
  1980 => x"849c80e9",
  1981 => x"51bad52d",
  1982 => x"80dda008",
  1983 => x"802e8d38",
  1984 => x"bbc82dff",
  1985 => x"135372c6",
  1986 => x"38bed504",
  1987 => x"81ff0bd4",
  1988 => x"0c80dda0",
  1989 => x"085287fc",
  1990 => x"80fa51ba",
  1991 => x"d52d80dd",
  1992 => x"a008b238",
  1993 => x"81ff0bd4",
  1994 => x"0cd40853",
  1995 => x"81ff0bd4",
  1996 => x"0c81ff0b",
  1997 => x"d40c81ff",
  1998 => x"0bd40c81",
  1999 => x"ff0bd40c",
  2000 => x"72862a70",
  2001 => x"81067656",
  2002 => x"51537296",
  2003 => x"3880dda0",
  2004 => x"0854bee2",
  2005 => x"0473822e",
  2006 => x"fedb38ff",
  2007 => x"145473fe",
  2008 => x"e7387380",
  2009 => x"de8c0c73",
  2010 => x"8b388152",
  2011 => x"87fc80d0",
  2012 => x"51bad52d",
  2013 => x"81ff0bd4",
  2014 => x"0cd00870",
  2015 => x"8f2a7081",
  2016 => x"06515153",
  2017 => x"72f33872",
  2018 => x"d00c81ff",
  2019 => x"0bd40c81",
  2020 => x"537280dd",
  2021 => x"a00c0294",
  2022 => x"050d0402",
  2023 => x"e8050d78",
  2024 => x"55805681",
  2025 => x"ff0bd40c",
  2026 => x"d008708f",
  2027 => x"2a708106",
  2028 => x"51515372",
  2029 => x"f3388281",
  2030 => x"0bd00c81",
  2031 => x"ff0bd40c",
  2032 => x"775287fc",
  2033 => x"80d151ba",
  2034 => x"d52d80db",
  2035 => x"c6df5480",
  2036 => x"dda00880",
  2037 => x"2e8c3880",
  2038 => x"d7f85186",
  2039 => x"a02d80c0",
  2040 => x"b70481ff",
  2041 => x"0bd40cd4",
  2042 => x"087081ff",
  2043 => x"06515372",
  2044 => x"81fe2e09",
  2045 => x"81069f38",
  2046 => x"80ff53ba",
  2047 => x"862d80dd",
  2048 => x"a0087570",
  2049 => x"8405570c",
  2050 => x"ff135372",
  2051 => x"8025ec38",
  2052 => x"815680c0",
  2053 => x"9c04ff14",
  2054 => x"5473c738",
  2055 => x"81ff0bd4",
  2056 => x"0c81ff0b",
  2057 => x"d40cd008",
  2058 => x"708f2a70",
  2059 => x"81065151",
  2060 => x"5372f338",
  2061 => x"72d00c75",
  2062 => x"80dda00c",
  2063 => x"0298050d",
  2064 => x"0402e805",
  2065 => x"0d77797b",
  2066 => x"58555580",
  2067 => x"53727625",
  2068 => x"a5387470",
  2069 => x"81055680",
  2070 => x"f52d7470",
  2071 => x"81055680",
  2072 => x"f52d5252",
  2073 => x"71712e87",
  2074 => x"38815180",
  2075 => x"c0f80481",
  2076 => x"135380c0",
  2077 => x"cd048051",
  2078 => x"7080dda0",
  2079 => x"0c029805",
  2080 => x"0d0402ec",
  2081 => x"050d7655",
  2082 => x"74802e80",
  2083 => x"c4389a15",
  2084 => x"80e02d51",
  2085 => x"80cfb62d",
  2086 => x"80dda008",
  2087 => x"80dda008",
  2088 => x"80e4c00c",
  2089 => x"80dda008",
  2090 => x"545480e4",
  2091 => x"9c08802e",
  2092 => x"9b389415",
  2093 => x"80e02d51",
  2094 => x"80cfb62d",
  2095 => x"80dda008",
  2096 => x"902b83ff",
  2097 => x"f00a0670",
  2098 => x"75075153",
  2099 => x"7280e4c0",
  2100 => x"0c80e4c0",
  2101 => x"08537280",
  2102 => x"2e9e3880",
  2103 => x"e49408fe",
  2104 => x"14712980",
  2105 => x"e4a80805",
  2106 => x"80e4c40c",
  2107 => x"70842b80",
  2108 => x"e4a00c54",
  2109 => x"80c2a704",
  2110 => x"80e4ac08",
  2111 => x"80e4c00c",
  2112 => x"80e4b008",
  2113 => x"80e4c40c",
  2114 => x"80e49c08",
  2115 => x"802e8c38",
  2116 => x"80e49408",
  2117 => x"842b5380",
  2118 => x"c2a20480",
  2119 => x"e4b40884",
  2120 => x"2b537280",
  2121 => x"e4a00c02",
  2122 => x"94050d04",
  2123 => x"02d8050d",
  2124 => x"800b80e4",
  2125 => x"9c0c8454",
  2126 => x"bc992d80",
  2127 => x"dda00880",
  2128 => x"2e983880",
  2129 => x"de905280",
  2130 => x"51bf9b2d",
  2131 => x"80dda008",
  2132 => x"802e8738",
  2133 => x"fe5480c2",
  2134 => x"e204ff14",
  2135 => x"54738024",
  2136 => x"d738738e",
  2137 => x"3880d888",
  2138 => x"5186a02d",
  2139 => x"735580c8",
  2140 => x"c5048056",
  2141 => x"810b80e4",
  2142 => x"c80c8853",
  2143 => x"80d89c52",
  2144 => x"80dec651",
  2145 => x"80c0c12d",
  2146 => x"80dda008",
  2147 => x"762e0981",
  2148 => x"06893880",
  2149 => x"dda00880",
  2150 => x"e4c80c88",
  2151 => x"5380d8a8",
  2152 => x"5280dee2",
  2153 => x"5180c0c1",
  2154 => x"2d80dda0",
  2155 => x"08893880",
  2156 => x"dda00880",
  2157 => x"e4c80c80",
  2158 => x"e4c80880",
  2159 => x"2e818438",
  2160 => x"80e1d60b",
  2161 => x"80f52d80",
  2162 => x"e1d70b80",
  2163 => x"f52d7198",
  2164 => x"2b71902b",
  2165 => x"0780e1d8",
  2166 => x"0b80f52d",
  2167 => x"70882b72",
  2168 => x"0780e1d9",
  2169 => x"0b80f52d",
  2170 => x"710780e2",
  2171 => x"8e0b80f5",
  2172 => x"2d80e28f",
  2173 => x"0b80f52d",
  2174 => x"71882b07",
  2175 => x"535f5452",
  2176 => x"5a565755",
  2177 => x"7381abaa",
  2178 => x"2e098106",
  2179 => x"90387551",
  2180 => x"80cf852d",
  2181 => x"80dda008",
  2182 => x"5680c4ac",
  2183 => x"047382d4",
  2184 => x"d52e8938",
  2185 => x"80d8b451",
  2186 => x"80c4fb04",
  2187 => x"80de9052",
  2188 => x"7551bf9b",
  2189 => x"2d80dda0",
  2190 => x"085580dd",
  2191 => x"a008802e",
  2192 => x"84833888",
  2193 => x"5380d8a8",
  2194 => x"5280dee2",
  2195 => x"5180c0c1",
  2196 => x"2d80dda0",
  2197 => x"088b3881",
  2198 => x"0b80e49c",
  2199 => x"0c80c582",
  2200 => x"04885380",
  2201 => x"d89c5280",
  2202 => x"dec65180",
  2203 => x"c0c12d80",
  2204 => x"dda00880",
  2205 => x"2e8c3880",
  2206 => x"d8c85186",
  2207 => x"a02d80c5",
  2208 => x"e10480e2",
  2209 => x"8e0b80f5",
  2210 => x"2d547380",
  2211 => x"d52e0981",
  2212 => x"0680ce38",
  2213 => x"80e28f0b",
  2214 => x"80f52d54",
  2215 => x"7381aa2e",
  2216 => x"098106bd",
  2217 => x"38800b80",
  2218 => x"de900b80",
  2219 => x"f52d5654",
  2220 => x"7481e92e",
  2221 => x"83388154",
  2222 => x"7481eb2e",
  2223 => x"8c388055",
  2224 => x"73752e09",
  2225 => x"810682fd",
  2226 => x"3880de9b",
  2227 => x"0b80f52d",
  2228 => x"55748e38",
  2229 => x"80de9c0b",
  2230 => x"80f52d54",
  2231 => x"73822e87",
  2232 => x"38805580",
  2233 => x"c8c50480",
  2234 => x"de9d0b80",
  2235 => x"f52d7080",
  2236 => x"e4940cff",
  2237 => x"0580e498",
  2238 => x"0c80de9e",
  2239 => x"0b80f52d",
  2240 => x"80de9f0b",
  2241 => x"80f52d58",
  2242 => x"76057782",
  2243 => x"80290570",
  2244 => x"80e4a40c",
  2245 => x"80dea00b",
  2246 => x"80f52d70",
  2247 => x"80e4b80c",
  2248 => x"80e49c08",
  2249 => x"59575876",
  2250 => x"802e81b9",
  2251 => x"38885380",
  2252 => x"d8a85280",
  2253 => x"dee25180",
  2254 => x"c0c12d80",
  2255 => x"dda00882",
  2256 => x"843880e4",
  2257 => x"94087084",
  2258 => x"2b80e4a0",
  2259 => x"0c7080e4",
  2260 => x"b40c80de",
  2261 => x"b50b80f5",
  2262 => x"2d80deb4",
  2263 => x"0b80f52d",
  2264 => x"71828029",
  2265 => x"0580deb6",
  2266 => x"0b80f52d",
  2267 => x"70848080",
  2268 => x"291280de",
  2269 => x"b70b80f5",
  2270 => x"2d708180",
  2271 => x"0a291270",
  2272 => x"80e4bc0c",
  2273 => x"80e4b808",
  2274 => x"712980e4",
  2275 => x"a4080570",
  2276 => x"80e4a80c",
  2277 => x"80debd0b",
  2278 => x"80f52d80",
  2279 => x"debc0b80",
  2280 => x"f52d7182",
  2281 => x"80290580",
  2282 => x"debe0b80",
  2283 => x"f52d7084",
  2284 => x"80802912",
  2285 => x"80debf0b",
  2286 => x"80f52d70",
  2287 => x"982b81f0",
  2288 => x"0a067205",
  2289 => x"7080e4ac",
  2290 => x"0cfe117e",
  2291 => x"29770580",
  2292 => x"e4b00c52",
  2293 => x"59524354",
  2294 => x"5e515259",
  2295 => x"525d5759",
  2296 => x"5780c8bd",
  2297 => x"0480dea2",
  2298 => x"0b80f52d",
  2299 => x"80dea10b",
  2300 => x"80f52d71",
  2301 => x"82802905",
  2302 => x"7080e4a0",
  2303 => x"0c70a029",
  2304 => x"83ff0570",
  2305 => x"892a7080",
  2306 => x"e4b40c80",
  2307 => x"dea70b80",
  2308 => x"f52d80de",
  2309 => x"a60b80f5",
  2310 => x"2d718280",
  2311 => x"29057080",
  2312 => x"e4bc0c7b",
  2313 => x"71291e70",
  2314 => x"80e4b00c",
  2315 => x"7d80e4ac",
  2316 => x"0c730580",
  2317 => x"e4a80c55",
  2318 => x"5e515155",
  2319 => x"55805180",
  2320 => x"c1822d81",
  2321 => x"557480dd",
  2322 => x"a00c02a8",
  2323 => x"050d0402",
  2324 => x"ec050d76",
  2325 => x"70872c71",
  2326 => x"80ff0655",
  2327 => x"565480e4",
  2328 => x"9c088a38",
  2329 => x"73882c74",
  2330 => x"81ff0654",
  2331 => x"5580de90",
  2332 => x"5280e4a4",
  2333 => x"081551bf",
  2334 => x"9b2d80dd",
  2335 => x"a0085480",
  2336 => x"dda00880",
  2337 => x"2ebb3880",
  2338 => x"e49c0880",
  2339 => x"2e9c3872",
  2340 => x"842980de",
  2341 => x"90057008",
  2342 => x"525380cf",
  2343 => x"852d80dd",
  2344 => x"a008f00a",
  2345 => x"065380c9",
  2346 => x"bf047210",
  2347 => x"80de9005",
  2348 => x"7080e02d",
  2349 => x"525380cf",
  2350 => x"b62d80dd",
  2351 => x"a0085372",
  2352 => x"547380dd",
  2353 => x"a00c0294",
  2354 => x"050d0402",
  2355 => x"e0050d79",
  2356 => x"70842c80",
  2357 => x"e4c40805",
  2358 => x"718f0652",
  2359 => x"5553728a",
  2360 => x"3880de90",
  2361 => x"527351bf",
  2362 => x"9b2d72a0",
  2363 => x"2980de90",
  2364 => x"05548074",
  2365 => x"80f52d56",
  2366 => x"5374732e",
  2367 => x"83388153",
  2368 => x"7481e52e",
  2369 => x"81f53881",
  2370 => x"70740654",
  2371 => x"5872802e",
  2372 => x"81e9388b",
  2373 => x"1480f52d",
  2374 => x"70832a79",
  2375 => x"06585676",
  2376 => x"9c3880db",
  2377 => x"e4085372",
  2378 => x"89387280",
  2379 => x"e2900b81",
  2380 => x"b72d7680",
  2381 => x"dbe40c73",
  2382 => x"5380cbfd",
  2383 => x"04758f2e",
  2384 => x"09810681",
  2385 => x"b638749f",
  2386 => x"068d2980",
  2387 => x"e2831151",
  2388 => x"53811480",
  2389 => x"f52d7370",
  2390 => x"81055581",
  2391 => x"b72d8314",
  2392 => x"80f52d73",
  2393 => x"70810555",
  2394 => x"81b72d85",
  2395 => x"1480f52d",
  2396 => x"73708105",
  2397 => x"5581b72d",
  2398 => x"871480f5",
  2399 => x"2d737081",
  2400 => x"055581b7",
  2401 => x"2d891480",
  2402 => x"f52d7370",
  2403 => x"81055581",
  2404 => x"b72d8e14",
  2405 => x"80f52d73",
  2406 => x"70810555",
  2407 => x"81b72d90",
  2408 => x"1480f52d",
  2409 => x"73708105",
  2410 => x"5581b72d",
  2411 => x"921480f5",
  2412 => x"2d737081",
  2413 => x"055581b7",
  2414 => x"2d941480",
  2415 => x"f52d7370",
  2416 => x"81055581",
  2417 => x"b72d9614",
  2418 => x"80f52d73",
  2419 => x"70810555",
  2420 => x"81b72d98",
  2421 => x"1480f52d",
  2422 => x"73708105",
  2423 => x"5581b72d",
  2424 => x"9c1480f5",
  2425 => x"2d737081",
  2426 => x"055581b7",
  2427 => x"2d9e1480",
  2428 => x"f52d7381",
  2429 => x"b72d7780",
  2430 => x"dbe40c80",
  2431 => x"537280dd",
  2432 => x"a00c02a0",
  2433 => x"050d0402",
  2434 => x"cc050d7e",
  2435 => x"605e5a80",
  2436 => x"0b80e4c0",
  2437 => x"0880e4c4",
  2438 => x"08595c56",
  2439 => x"805880e4",
  2440 => x"a008782e",
  2441 => x"81bd3877",
  2442 => x"8f06a017",
  2443 => x"57547391",
  2444 => x"3880de90",
  2445 => x"52765181",
  2446 => x"1757bf9b",
  2447 => x"2d80de90",
  2448 => x"56807680",
  2449 => x"f52d5654",
  2450 => x"74742e83",
  2451 => x"38815474",
  2452 => x"81e52e81",
  2453 => x"82388170",
  2454 => x"7506555c",
  2455 => x"73802e80",
  2456 => x"f6388b16",
  2457 => x"80f52d98",
  2458 => x"06597880",
  2459 => x"ea388b53",
  2460 => x"7c527551",
  2461 => x"80c0c12d",
  2462 => x"80dda008",
  2463 => x"80d9389c",
  2464 => x"16085180",
  2465 => x"cf852d80",
  2466 => x"dda00884",
  2467 => x"1b0c9a16",
  2468 => x"80e02d51",
  2469 => x"80cfb62d",
  2470 => x"80dda008",
  2471 => x"80dda008",
  2472 => x"881c0c80",
  2473 => x"dda00855",
  2474 => x"5580e49c",
  2475 => x"08802e9a",
  2476 => x"38941680",
  2477 => x"e02d5180",
  2478 => x"cfb62d80",
  2479 => x"dda00890",
  2480 => x"2b83fff0",
  2481 => x"0a067016",
  2482 => x"51547388",
  2483 => x"1b0c787a",
  2484 => x"0c7b5480",
  2485 => x"cea10481",
  2486 => x"185880e4",
  2487 => x"a0087826",
  2488 => x"fec53880",
  2489 => x"e49c0880",
  2490 => x"2eb5387a",
  2491 => x"5180c8cf",
  2492 => x"2d80dda0",
  2493 => x"0880dda0",
  2494 => x"0880ffff",
  2495 => x"fff80655",
  2496 => x"5b7380ff",
  2497 => x"fffff82e",
  2498 => x"963880dd",
  2499 => x"a008fe05",
  2500 => x"80e49408",
  2501 => x"2980e4a8",
  2502 => x"08055780",
  2503 => x"cc9c0480",
  2504 => x"547380dd",
  2505 => x"a00c02b4",
  2506 => x"050d0402",
  2507 => x"f4050d74",
  2508 => x"70088105",
  2509 => x"710c7008",
  2510 => x"80e49808",
  2511 => x"06535371",
  2512 => x"90388813",
  2513 => x"085180c8",
  2514 => x"cf2d80dd",
  2515 => x"a0088814",
  2516 => x"0c810b80",
  2517 => x"dda00c02",
  2518 => x"8c050d04",
  2519 => x"02f0050d",
  2520 => x"75881108",
  2521 => x"fe0580e4",
  2522 => x"94082980",
  2523 => x"e4a80811",
  2524 => x"720880e4",
  2525 => x"98080605",
  2526 => x"79555354",
  2527 => x"54bf9b2d",
  2528 => x"0290050d",
  2529 => x"0402f405",
  2530 => x"0d747088",
  2531 => x"2a83fe80",
  2532 => x"06707298",
  2533 => x"2a077288",
  2534 => x"2b87fc80",
  2535 => x"80067398",
  2536 => x"2b81f00a",
  2537 => x"06717307",
  2538 => x"0780dda0",
  2539 => x"0c565153",
  2540 => x"51028c05",
  2541 => x"0d0402f8",
  2542 => x"050d028e",
  2543 => x"0580f52d",
  2544 => x"74882b07",
  2545 => x"7083ffff",
  2546 => x"0680dda0",
  2547 => x"0c510288",
  2548 => x"050d0402",
  2549 => x"f4050d74",
  2550 => x"76785354",
  2551 => x"52807125",
  2552 => x"97387270",
  2553 => x"81055480",
  2554 => x"f52d7270",
  2555 => x"81055481",
  2556 => x"b72dff11",
  2557 => x"5170eb38",
  2558 => x"807281b7",
  2559 => x"2d028c05",
  2560 => x"0d0402e8",
  2561 => x"050d7756",
  2562 => x"80705654",
  2563 => x"737624b7",
  2564 => x"3880e4a0",
  2565 => x"08742eaf",
  2566 => x"38735180",
  2567 => x"c9cb2d80",
  2568 => x"dda00880",
  2569 => x"dda00809",
  2570 => x"81057080",
  2571 => x"dda00807",
  2572 => x"9f2a7705",
  2573 => x"81175757",
  2574 => x"53537476",
  2575 => x"24893880",
  2576 => x"e4a00874",
  2577 => x"26d33872",
  2578 => x"80dda00c",
  2579 => x"0298050d",
  2580 => x"0402f005",
  2581 => x"0d80dd9c",
  2582 => x"08165180",
  2583 => x"d0822d80",
  2584 => x"dda00880",
  2585 => x"2ea0388b",
  2586 => x"5380dda0",
  2587 => x"085280e2",
  2588 => x"905180cf",
  2589 => x"d32d80e4",
  2590 => x"cc085473",
  2591 => x"802e8738",
  2592 => x"80e29051",
  2593 => x"732d0290",
  2594 => x"050d0402",
  2595 => x"dc050d80",
  2596 => x"705a5574",
  2597 => x"80dd9c08",
  2598 => x"25b53880",
  2599 => x"e4a00875",
  2600 => x"2ead3878",
  2601 => x"5180c9cb",
  2602 => x"2d80dda0",
  2603 => x"08098105",
  2604 => x"7080dda0",
  2605 => x"08079f2a",
  2606 => x"7605811b",
  2607 => x"5b565474",
  2608 => x"80dd9c08",
  2609 => x"25893880",
  2610 => x"e4a00879",
  2611 => x"26d53880",
  2612 => x"557880e4",
  2613 => x"a0082781",
  2614 => x"e4387851",
  2615 => x"80c9cb2d",
  2616 => x"80dda008",
  2617 => x"802e81b4",
  2618 => x"3880dda0",
  2619 => x"088b0580",
  2620 => x"f52d7084",
  2621 => x"2a708106",
  2622 => x"77107884",
  2623 => x"2b80e290",
  2624 => x"0b80f52d",
  2625 => x"5c5c5351",
  2626 => x"55567380",
  2627 => x"2e80ce38",
  2628 => x"7416822b",
  2629 => x"80d3e10b",
  2630 => x"80dbf012",
  2631 => x"0c547775",
  2632 => x"311080e4",
  2633 => x"d0115556",
  2634 => x"90747081",
  2635 => x"055681b7",
  2636 => x"2da07481",
  2637 => x"b72d7681",
  2638 => x"ff068116",
  2639 => x"58547380",
  2640 => x"2e8b389c",
  2641 => x"5380e290",
  2642 => x"5280d2d4",
  2643 => x"048b5380",
  2644 => x"dda00852",
  2645 => x"80e4d216",
  2646 => x"5180d392",
  2647 => x"04741682",
  2648 => x"2b80d0d1",
  2649 => x"0b80dbf0",
  2650 => x"120c5476",
  2651 => x"81ff0681",
  2652 => x"16585473",
  2653 => x"802e8b38",
  2654 => x"9c5380e2",
  2655 => x"905280d3",
  2656 => x"89048b53",
  2657 => x"80dda008",
  2658 => x"52777531",
  2659 => x"1080e4d0",
  2660 => x"05517655",
  2661 => x"80cfd32d",
  2662 => x"80d3b104",
  2663 => x"74902975",
  2664 => x"31701080",
  2665 => x"e4d00551",
  2666 => x"5480dda0",
  2667 => x"087481b7",
  2668 => x"2d811959",
  2669 => x"748b24a4",
  2670 => x"3880d1d1",
  2671 => x"04749029",
  2672 => x"75317010",
  2673 => x"80e4d005",
  2674 => x"8c773157",
  2675 => x"51548074",
  2676 => x"81b72d9e",
  2677 => x"14ff1656",
  2678 => x"5474f338",
  2679 => x"02a4050d",
  2680 => x"0402fc05",
  2681 => x"0d80dd9c",
  2682 => x"08135180",
  2683 => x"d0822d80",
  2684 => x"dda00880",
  2685 => x"2e8a3880",
  2686 => x"dda00851",
  2687 => x"80c1822d",
  2688 => x"800b80dd",
  2689 => x"9c0c80d1",
  2690 => x"8b2daf88",
  2691 => x"2d028405",
  2692 => x"0d0402fc",
  2693 => x"050d7251",
  2694 => x"70fd2eb2",
  2695 => x"3870fd24",
  2696 => x"8b3870fc",
  2697 => x"2e80d038",
  2698 => x"80d58104",
  2699 => x"70fe2eb9",
  2700 => x"3870ff2e",
  2701 => x"09810680",
  2702 => x"c83880dd",
  2703 => x"9c085170",
  2704 => x"802ebe38",
  2705 => x"ff1180dd",
  2706 => x"9c0c80d5",
  2707 => x"810480dd",
  2708 => x"9c08f405",
  2709 => x"7080dd9c",
  2710 => x"0c517080",
  2711 => x"25a33880",
  2712 => x"0b80dd9c",
  2713 => x"0c80d581",
  2714 => x"0480dd9c",
  2715 => x"08810580",
  2716 => x"dd9c0c80",
  2717 => x"d5810480",
  2718 => x"dd9c088c",
  2719 => x"0580dd9c",
  2720 => x"0c80d18b",
  2721 => x"2daf882d",
  2722 => x"0284050d",
  2723 => x"0402fc05",
  2724 => x"0d800b80",
  2725 => x"dd9c0c80",
  2726 => x"d18b2dae",
  2727 => x"842d80dd",
  2728 => x"a00880dd",
  2729 => x"8c0c80db",
  2730 => x"e851b0ae",
  2731 => x"2d028405",
  2732 => x"0d047180",
  2733 => x"e4cc0c04",
  2734 => x"00ffffff",
  2735 => x"ff00ffff",
  2736 => x"ffff00ff",
  2737 => x"ffffff00",
  2738 => x"30313233",
  2739 => x"34353637",
  2740 => x"38394142",
  2741 => x"43444546",
  2742 => x"00000000",
  2743 => x"52657365",
  2744 => x"74000000",
  2745 => x"5363616e",
  2746 => x"6c696e65",
  2747 => x"73000000",
  2748 => x"50414c20",
  2749 => x"2f204e54",
  2750 => x"53430000",
  2751 => x"436f6c6f",
  2752 => x"72000000",
  2753 => x"44696666",
  2754 => x"6963756c",
  2755 => x"74792041",
  2756 => x"00000000",
  2757 => x"44696666",
  2758 => x"6963756c",
  2759 => x"74792042",
  2760 => x"00000000",
  2761 => x"2a537570",
  2762 => x"65726368",
  2763 => x"69702069",
  2764 => x"6e206361",
  2765 => x"72747269",
  2766 => x"64676500",
  2767 => x"2a42616e",
  2768 => x"6b204530",
  2769 => x"00000000",
  2770 => x"2a42616e",
  2771 => x"6b204537",
  2772 => x"00000000",
  2773 => x"53656c65",
  2774 => x"63740000",
  2775 => x"53746172",
  2776 => x"74000000",
  2777 => x"4c6f6164",
  2778 => x"20524f4d",
  2779 => x"20100000",
  2780 => x"45786974",
  2781 => x"00000000",
  2782 => x"524f4d20",
  2783 => x"6c6f6164",
  2784 => x"696e6720",
  2785 => x"6661696c",
  2786 => x"65640000",
  2787 => x"4f4b0000",
  2788 => x"496e6974",
  2789 => x"69616c69",
  2790 => x"7a696e67",
  2791 => x"20534420",
  2792 => x"63617264",
  2793 => x"0a000000",
  2794 => x"16200000",
  2795 => x"14200000",
  2796 => x"15200000",
  2797 => x"53442069",
  2798 => x"6e69742e",
  2799 => x"2e2e0a00",
  2800 => x"53442063",
  2801 => x"61726420",
  2802 => x"72657365",
  2803 => x"74206661",
  2804 => x"696c6564",
  2805 => x"210a0000",
  2806 => x"53444843",
  2807 => x"20657272",
  2808 => x"6f72210a",
  2809 => x"00000000",
  2810 => x"57726974",
  2811 => x"65206661",
  2812 => x"696c6564",
  2813 => x"0a000000",
  2814 => x"52656164",
  2815 => x"20666169",
  2816 => x"6c65640a",
  2817 => x"00000000",
  2818 => x"43617264",
  2819 => x"20696e69",
  2820 => x"74206661",
  2821 => x"696c6564",
  2822 => x"0a000000",
  2823 => x"46415431",
  2824 => x"36202020",
  2825 => x"00000000",
  2826 => x"46415433",
  2827 => x"32202020",
  2828 => x"00000000",
  2829 => x"4e6f2070",
  2830 => x"61727469",
  2831 => x"74696f6e",
  2832 => x"20736967",
  2833 => x"0a000000",
  2834 => x"42616420",
  2835 => x"70617274",
  2836 => x"0a000000",
  2837 => x"4261636b",
  2838 => x"00000000",
  2839 => x"00000002",
  2840 => x"00000002",
  2841 => x"00002adc",
  2842 => x"0000035a",
  2843 => x"00000001",
  2844 => x"00002ae4",
  2845 => x"00000000",
  2846 => x"00000001",
  2847 => x"00002af0",
  2848 => x"00000001",
  2849 => x"00000001",
  2850 => x"00002afc",
  2851 => x"00000002",
  2852 => x"00000001",
  2853 => x"00002b04",
  2854 => x"00000003",
  2855 => x"00000001",
  2856 => x"00002b14",
  2857 => x"00000004",
  2858 => x"00000001",
  2859 => x"00002b24",
  2860 => x"00000005",
  2861 => x"00000001",
  2862 => x"00002b3c",
  2863 => x"00000008",
  2864 => x"00000001",
  2865 => x"00002b48",
  2866 => x"00000009",
  2867 => x"00000002",
  2868 => x"00002b54",
  2869 => x"0000036e",
  2870 => x"00000002",
  2871 => x"00002b5c",
  2872 => x"00000a3f",
  2873 => x"00000002",
  2874 => x"00002b64",
  2875 => x"00002a8d",
  2876 => x"00000002",
  2877 => x"00002b70",
  2878 => x"00001721",
  2879 => x"00000000",
  2880 => x"00000000",
  2881 => x"00000000",
  2882 => x"00000004",
  2883 => x"00002b78",
  2884 => x"00002d08",
  2885 => x"00000004",
  2886 => x"00002b8c",
  2887 => x"00002c60",
  2888 => x"00000000",
  2889 => x"00000000",
  2890 => x"00000000",
  2891 => x"00000000",
  2892 => x"00000000",
  2893 => x"00000000",
  2894 => x"00000000",
  2895 => x"00000000",
  2896 => x"00000000",
  2897 => x"00000000",
  2898 => x"00000000",
  2899 => x"00000000",
  2900 => x"00000000",
  2901 => x"00000000",
  2902 => x"00000000",
  2903 => x"00000000",
  2904 => x"00000000",
  2905 => x"00000000",
  2906 => x"00000000",
  2907 => x"761c1c1c",
  2908 => x"1c1c051c",
  2909 => x"1c1c1c1c",
  2910 => x"f2f5fafd",
  2911 => x"5a000000",
  2912 => x"00000000",
  2913 => x"00000000",
  2914 => x"00000000",
  2915 => x"00000000",
  2916 => x"00000000",
  2917 => x"00000000",
  2918 => x"00000000",
  2919 => x"00000000",
  2920 => x"00000000",
  2921 => x"00000000",
  2922 => x"00000000",
  2923 => x"00000000",
  2924 => x"00000000",
  2925 => x"00000000",
  2926 => x"00000000",
  2927 => x"00000000",
  2928 => x"00000000",
  2929 => x"00000000",
  2930 => x"0001ffff",
  2931 => x"0001ffff",
  2932 => x"0001ffff",
  2933 => x"00000000",
  2934 => x"00000000",
  2935 => x"00000006",
  2936 => x"00000000",
  2937 => x"00000000",
  2938 => x"00000002",
  2939 => x"00003250",
  2940 => x"00002851",
  2941 => x"00000002",
  2942 => x"0000326e",
  2943 => x"00002851",
  2944 => x"00000002",
  2945 => x"0000328c",
  2946 => x"00002851",
  2947 => x"00000002",
  2948 => x"000032aa",
  2949 => x"00002851",
  2950 => x"00000002",
  2951 => x"000032c8",
  2952 => x"00002851",
  2953 => x"00000002",
  2954 => x"000032e6",
  2955 => x"00002851",
  2956 => x"00000002",
  2957 => x"00003304",
  2958 => x"00002851",
  2959 => x"00000002",
  2960 => x"00003322",
  2961 => x"00002851",
  2962 => x"00000002",
  2963 => x"00003340",
  2964 => x"00002851",
  2965 => x"00000002",
  2966 => x"0000335e",
  2967 => x"00002851",
  2968 => x"00000002",
  2969 => x"0000337c",
  2970 => x"00002851",
  2971 => x"00000002",
  2972 => x"0000339a",
  2973 => x"00002851",
  2974 => x"00000002",
  2975 => x"000033b8",
  2976 => x"00002851",
  2977 => x"00000004",
  2978 => x"00002c54",
  2979 => x"00000000",
  2980 => x"00000000",
  2981 => x"00000000",
  2982 => x"00002a12",
  2983 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

