-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80dc",
     9 => x"90080b0b",
    10 => x"80dc9408",
    11 => x"0b0b80dc",
    12 => x"98080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"dc980c0b",
    16 => x"0b80dc94",
    17 => x"0c0b0b80",
    18 => x"dc900c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d4d4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80dc9070",
    57 => x"80e7d027",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a5ed",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80dc",
    65 => x"a00c9f0b",
    66 => x"80dca40c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"dca408ff",
    70 => x"0580dca4",
    71 => x"0c80dca4",
    72 => x"088025e8",
    73 => x"3880dca0",
    74 => x"08ff0580",
    75 => x"dca00c80",
    76 => x"dca00880",
    77 => x"25d03880",
    78 => x"0b80dca4",
    79 => x"0c800b80",
    80 => x"dca00c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80dca008",
   100 => x"25913882",
   101 => x"c82d80dc",
   102 => x"a008ff05",
   103 => x"80dca00c",
   104 => x"838a0480",
   105 => x"dca00880",
   106 => x"dca40853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80dca008",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"dca40881",
   116 => x"0580dca4",
   117 => x"0c80dca4",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80dca4",
   121 => x"0c80dca0",
   122 => x"08810580",
   123 => x"dca00c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480dc",
   128 => x"a4088105",
   129 => x"80dca40c",
   130 => x"80dca408",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80dca4",
   134 => x"0c80dca0",
   135 => x"08810580",
   136 => x"dca00c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"dca80cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"dca80c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280dc",
   177 => x"a8088407",
   178 => x"80dca80c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80d8",
   183 => x"840c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80dca8",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80dc",
   208 => x"900c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02f8050d",
  1093 => x"028f0580",
  1094 => x"f52d80d8",
  1095 => x"8c085252",
  1096 => x"7080ddbd",
  1097 => x"279a3871",
  1098 => x"7181b72d",
  1099 => x"80d88c08",
  1100 => x"810580d8",
  1101 => x"8c0c80d8",
  1102 => x"8c085180",
  1103 => x"7181b72d",
  1104 => x"0288050d",
  1105 => x"0402f405",
  1106 => x"0d747084",
  1107 => x"2a708f06",
  1108 => x"80d88808",
  1109 => x"057080f5",
  1110 => x"2d545153",
  1111 => x"53a2902d",
  1112 => x"728f0680",
  1113 => x"d8880805",
  1114 => x"7080f52d",
  1115 => x"5253a290",
  1116 => x"2d028c05",
  1117 => x"0d0402f4",
  1118 => x"050d7476",
  1119 => x"54527270",
  1120 => x"81055480",
  1121 => x"f52d5170",
  1122 => x"72708105",
  1123 => x"5481b72d",
  1124 => x"70ec3870",
  1125 => x"7281b72d",
  1126 => x"028c050d",
  1127 => x"0402d005",
  1128 => x"0d800b80",
  1129 => x"dacc0881",
  1130 => x"8006715d",
  1131 => x"5d59810b",
  1132 => x"ec0c840b",
  1133 => x"ec0c7d52",
  1134 => x"80dcac51",
  1135 => x"80cba32d",
  1136 => x"80dc9008",
  1137 => x"792e80ff",
  1138 => x"3880dcb0",
  1139 => x"0879ff12",
  1140 => x"57595774",
  1141 => x"792e8b38",
  1142 => x"81187581",
  1143 => x"2a565874",
  1144 => x"f738f718",
  1145 => x"58815980",
  1146 => x"772580db",
  1147 => x"38775274",
  1148 => x"5184a82d",
  1149 => x"80de8852",
  1150 => x"80dcac51",
  1151 => x"80cdf72d",
  1152 => x"80dc9008",
  1153 => x"802ea638",
  1154 => x"80de885a",
  1155 => x"7ba73883",
  1156 => x"ff567970",
  1157 => x"81055b80",
  1158 => x"f52d7b81",
  1159 => x"1d5de40c",
  1160 => x"e80cff16",
  1161 => x"56758025",
  1162 => x"e938a4b5",
  1163 => x"0480dc90",
  1164 => x"08598480",
  1165 => x"5780dcac",
  1166 => x"5180cdc6",
  1167 => x"2dfc8017",
  1168 => x"81165657",
  1169 => x"a3e70480",
  1170 => x"dcb008f8",
  1171 => x"0c810be0",
  1172 => x"0c805186",
  1173 => x"da2d86c7",
  1174 => x"2d78802e",
  1175 => x"883880d8",
  1176 => x"9051a4e9",
  1177 => x"0480d9c4",
  1178 => x"51afd22d",
  1179 => x"7880dc90",
  1180 => x"0c02b005",
  1181 => x"0d0402ec",
  1182 => x"050d80dc",
  1183 => x"fc0b80d8",
  1184 => x"8c0c80dc",
  1185 => x"fc538073",
  1186 => x"81b72d80",
  1187 => x"d9e80851",
  1188 => x"a2c52dba",
  1189 => x"51a2902d",
  1190 => x"ffb408ff",
  1191 => x"b8087098",
  1192 => x"2a535155",
  1193 => x"a2c52d74",
  1194 => x"902a7081",
  1195 => x"ff065254",
  1196 => x"a2c52d74",
  1197 => x"882a7081",
  1198 => x"ff065254",
  1199 => x"a2c52d74",
  1200 => x"81ff0651",
  1201 => x"a2c52d72",
  1202 => x"5280dcb8",
  1203 => x"51a2f62d",
  1204 => x"80d89051",
  1205 => x"afd22d80",
  1206 => x"d9e80884",
  1207 => x"0580d9e8",
  1208 => x"0c029405",
  1209 => x"0d04800b",
  1210 => x"80d9e80c",
  1211 => x"0402ec05",
  1212 => x"0d840bec",
  1213 => x"0cad8f2d",
  1214 => x"a7f52d81",
  1215 => x"f92d8353",
  1216 => x"acf22d81",
  1217 => x"51858d2d",
  1218 => x"ff135372",
  1219 => x"8025f138",
  1220 => x"840bec0c",
  1221 => x"80d6a851",
  1222 => x"86a02d80",
  1223 => x"c1cd2d80",
  1224 => x"dc900880",
  1225 => x"2e81b738",
  1226 => x"a39d5180",
  1227 => x"d4cd2d80",
  1228 => x"d6c05280",
  1229 => x"dcb851a2",
  1230 => x"f62d80d8",
  1231 => x"9051afd2",
  1232 => x"2dadb12d",
  1233 => x"a8c62daf",
  1234 => x"e52d80d8",
  1235 => x"a40b80f5",
  1236 => x"2d80dacc",
  1237 => x"08708106",
  1238 => x"55565472",
  1239 => x"802e8538",
  1240 => x"73840754",
  1241 => x"74812a70",
  1242 => x"81065153",
  1243 => x"72802e85",
  1244 => x"38738207",
  1245 => x"5474822a",
  1246 => x"70810651",
  1247 => x"5372802e",
  1248 => x"85387381",
  1249 => x"07547483",
  1250 => x"2a708106",
  1251 => x"51537280",
  1252 => x"2e853873",
  1253 => x"88075474",
  1254 => x"842a7081",
  1255 => x"06515372",
  1256 => x"802e8538",
  1257 => x"73900754",
  1258 => x"74852a70",
  1259 => x"81065153",
  1260 => x"72802e85",
  1261 => x"3873a007",
  1262 => x"5474882a",
  1263 => x"70810651",
  1264 => x"5372802e",
  1265 => x"86387380",
  1266 => x"c0075473",
  1267 => x"fc0c8653",
  1268 => x"80dc9008",
  1269 => x"83388453",
  1270 => x"72ec0ca6",
  1271 => x"c404800b",
  1272 => x"80dc900c",
  1273 => x"0294050d",
  1274 => x"0471980c",
  1275 => x"04ffb008",
  1276 => x"80dc900c",
  1277 => x"04810bff",
  1278 => x"b00c0480",
  1279 => x"0bffb00c",
  1280 => x"0402f805",
  1281 => x"0dffb408",
  1282 => x"709fff06",
  1283 => x"51517080",
  1284 => x"dabc082e",
  1285 => x"8c387080",
  1286 => x"dabc0c80",
  1287 => x"0b80dab8",
  1288 => x"0c80dab8",
  1289 => x"08518152",
  1290 => x"7087e82e",
  1291 => x"8f387087",
  1292 => x"e8248738",
  1293 => x"711180da",
  1294 => x"b80c8052",
  1295 => x"7180dc90",
  1296 => x"0c028805",
  1297 => x"0d0402e0",
  1298 => x"050da9d4",
  1299 => x"0480dc90",
  1300 => x"0881f02e",
  1301 => x"0981068a",
  1302 => x"38810b80",
  1303 => x"dac40ca9",
  1304 => x"d40480dc",
  1305 => x"900881e0",
  1306 => x"2e098106",
  1307 => x"8a38810b",
  1308 => x"80dac80c",
  1309 => x"a9d40480",
  1310 => x"dc900852",
  1311 => x"80dac808",
  1312 => x"802e8938",
  1313 => x"80dc9008",
  1314 => x"81800552",
  1315 => x"71842c72",
  1316 => x"8f065353",
  1317 => x"80dac408",
  1318 => x"802e9a38",
  1319 => x"72842980",
  1320 => x"d9ec0572",
  1321 => x"1381712b",
  1322 => x"70097308",
  1323 => x"06730c51",
  1324 => x"5353a9c8",
  1325 => x"04728429",
  1326 => x"80d9ec05",
  1327 => x"72138371",
  1328 => x"2b720807",
  1329 => x"720c5353",
  1330 => x"800b80da",
  1331 => x"c80c800b",
  1332 => x"80dac40c",
  1333 => x"80ddc051",
  1334 => x"abe52d80",
  1335 => x"dc9008ff",
  1336 => x"24feea38",
  1337 => x"a8812d80",
  1338 => x"dc900880",
  1339 => x"2e80ff38",
  1340 => x"8156800b",
  1341 => x"80dac008",
  1342 => x"80dabc08",
  1343 => x"80dac408",
  1344 => x"57595955",
  1345 => x"77760677",
  1346 => x"77065452",
  1347 => x"71732e80",
  1348 => x"c4387280",
  1349 => x"daac1680",
  1350 => x"f52d7084",
  1351 => x"2c718f06",
  1352 => x"52555354",
  1353 => x"73802e9a",
  1354 => x"38728429",
  1355 => x"80d9ec05",
  1356 => x"72138171",
  1357 => x"2b700973",
  1358 => x"0806730c",
  1359 => x"515353aa",
  1360 => x"d5047284",
  1361 => x"2980d9ec",
  1362 => x"05721383",
  1363 => x"712b7208",
  1364 => x"07720c53",
  1365 => x"53751081",
  1366 => x"1656568b",
  1367 => x"7525ffa4",
  1368 => x"387380da",
  1369 => x"c40c80da",
  1370 => x"bc0880da",
  1371 => x"c00c800b",
  1372 => x"80dc900c",
  1373 => x"02a0050d",
  1374 => x"0402f805",
  1375 => x"0d80d9ec",
  1376 => x"528f5180",
  1377 => x"72708405",
  1378 => x"540cff11",
  1379 => x"51708025",
  1380 => x"f2380288",
  1381 => x"050d0402",
  1382 => x"f0050d75",
  1383 => x"51a7fb2d",
  1384 => x"70822cfc",
  1385 => x"0680d9ec",
  1386 => x"1172109e",
  1387 => x"06710870",
  1388 => x"722a7083",
  1389 => x"0682742b",
  1390 => x"70097406",
  1391 => x"760c5451",
  1392 => x"56575351",
  1393 => x"53a7f52d",
  1394 => x"7180dc90",
  1395 => x"0c029005",
  1396 => x"0d0402fc",
  1397 => x"050d7251",
  1398 => x"80710c80",
  1399 => x"0b84120c",
  1400 => x"0284050d",
  1401 => x"0402f005",
  1402 => x"0d757008",
  1403 => x"84120853",
  1404 => x"5353ff54",
  1405 => x"71712ea8",
  1406 => x"38a7fb2d",
  1407 => x"84130870",
  1408 => x"84291488",
  1409 => x"11700870",
  1410 => x"81ff0684",
  1411 => x"18088111",
  1412 => x"8706841a",
  1413 => x"0c535155",
  1414 => x"515151a7",
  1415 => x"f52d7154",
  1416 => x"7380dc90",
  1417 => x"0c029005",
  1418 => x"0d0402f8",
  1419 => x"050da7fb",
  1420 => x"2de00870",
  1421 => x"8b2a7081",
  1422 => x"06515252",
  1423 => x"70802ea1",
  1424 => x"3880ddc0",
  1425 => x"08708429",
  1426 => x"80ddc805",
  1427 => x"7381ff06",
  1428 => x"710c5151",
  1429 => x"80ddc008",
  1430 => x"81118706",
  1431 => x"80ddc00c",
  1432 => x"51800b80",
  1433 => x"dde80ca7",
  1434 => x"ed2da7f5",
  1435 => x"2d028805",
  1436 => x"0d0402fc",
  1437 => x"050da7fb",
  1438 => x"2d810b80",
  1439 => x"dde80ca7",
  1440 => x"f52d80dd",
  1441 => x"e8085170",
  1442 => x"f9380284",
  1443 => x"050d0402",
  1444 => x"fc050d80",
  1445 => x"ddc051ab",
  1446 => x"d22daaf9",
  1447 => x"2dacaa51",
  1448 => x"a7e92d02",
  1449 => x"84050d04",
  1450 => x"80ddf408",
  1451 => x"80dc900c",
  1452 => x"0402fc05",
  1453 => x"0d810b80",
  1454 => x"dad00c81",
  1455 => x"51858d2d",
  1456 => x"0284050d",
  1457 => x"0402fc05",
  1458 => x"0dadcf04",
  1459 => x"a8c62d80",
  1460 => x"f651ab97",
  1461 => x"2d80dc90",
  1462 => x"08f23880",
  1463 => x"da51ab97",
  1464 => x"2d80dc90",
  1465 => x"08e63880",
  1466 => x"dc900880",
  1467 => x"dad00c80",
  1468 => x"dc900851",
  1469 => x"858d2d02",
  1470 => x"84050d04",
  1471 => x"02ec050d",
  1472 => x"76548052",
  1473 => x"870b8815",
  1474 => x"80f52d56",
  1475 => x"53747224",
  1476 => x"8338a053",
  1477 => x"72518384",
  1478 => x"2d81128b",
  1479 => x"1580f52d",
  1480 => x"54527272",
  1481 => x"25de3802",
  1482 => x"94050d04",
  1483 => x"02f0050d",
  1484 => x"80ddf408",
  1485 => x"5481f92d",
  1486 => x"800b80dd",
  1487 => x"f80c7308",
  1488 => x"802e8189",
  1489 => x"38820b80",
  1490 => x"dca40c80",
  1491 => x"ddf8088f",
  1492 => x"0680dca0",
  1493 => x"0c730852",
  1494 => x"71832e96",
  1495 => x"38718326",
  1496 => x"89387181",
  1497 => x"2eb038af",
  1498 => x"b6047185",
  1499 => x"2ea038af",
  1500 => x"b6048814",
  1501 => x"80f52d84",
  1502 => x"150880d6",
  1503 => x"d0535452",
  1504 => x"86a02d71",
  1505 => x"84291370",
  1506 => x"085252af",
  1507 => x"ba047351",
  1508 => x"adfc2daf",
  1509 => x"b60480da",
  1510 => x"cc088815",
  1511 => x"082c7081",
  1512 => x"06515271",
  1513 => x"802e8838",
  1514 => x"80d6d451",
  1515 => x"afb30480",
  1516 => x"d6d85186",
  1517 => x"a02d8414",
  1518 => x"085186a0",
  1519 => x"2d80ddf8",
  1520 => x"08810580",
  1521 => x"ddf80c8c",
  1522 => x"1454aebe",
  1523 => x"04029005",
  1524 => x"0d047180",
  1525 => x"ddf40cae",
  1526 => x"ac2d80dd",
  1527 => x"f808ff05",
  1528 => x"80ddfc0c",
  1529 => x"0402e805",
  1530 => x"0d80ddf4",
  1531 => x"0880de80",
  1532 => x"08575580",
  1533 => x"f651ab97",
  1534 => x"2d80dc90",
  1535 => x"08812a70",
  1536 => x"81065152",
  1537 => x"71802ea4",
  1538 => x"38b08f04",
  1539 => x"a8c62d80",
  1540 => x"f651ab97",
  1541 => x"2d80dc90",
  1542 => x"08f23880",
  1543 => x"dad00881",
  1544 => x"327080da",
  1545 => x"d00c7052",
  1546 => x"52858d2d",
  1547 => x"800b80dd",
  1548 => x"ec0c800b",
  1549 => x"80ddf00c",
  1550 => x"80dad008",
  1551 => x"838d3880",
  1552 => x"da51ab97",
  1553 => x"2d80dc90",
  1554 => x"08802e8c",
  1555 => x"3880ddec",
  1556 => x"08818007",
  1557 => x"80ddec0c",
  1558 => x"80d951ab",
  1559 => x"972d80dc",
  1560 => x"9008802e",
  1561 => x"8c3880dd",
  1562 => x"ec0880c0",
  1563 => x"0780ddec",
  1564 => x"0c819451",
  1565 => x"ab972d80",
  1566 => x"dc900880",
  1567 => x"2e8b3880",
  1568 => x"ddec0890",
  1569 => x"0780ddec",
  1570 => x"0c819151",
  1571 => x"ab972d80",
  1572 => x"dc900880",
  1573 => x"2e8b3880",
  1574 => x"ddec08a0",
  1575 => x"0780ddec",
  1576 => x"0c81f551",
  1577 => x"ab972d80",
  1578 => x"dc900880",
  1579 => x"2e8b3880",
  1580 => x"ddec0881",
  1581 => x"0780ddec",
  1582 => x"0c81f251",
  1583 => x"ab972d80",
  1584 => x"dc900880",
  1585 => x"2e8b3880",
  1586 => x"ddec0882",
  1587 => x"0780ddec",
  1588 => x"0c81eb51",
  1589 => x"ab972d80",
  1590 => x"dc900880",
  1591 => x"2e8b3880",
  1592 => x"ddec0884",
  1593 => x"0780ddec",
  1594 => x"0c81f451",
  1595 => x"ab972d80",
  1596 => x"dc900880",
  1597 => x"2e8b3880",
  1598 => x"ddec0888",
  1599 => x"0780ddec",
  1600 => x"0c80d851",
  1601 => x"ab972d80",
  1602 => x"dc900880",
  1603 => x"2e8c3880",
  1604 => x"ddf00881",
  1605 => x"800780dd",
  1606 => x"f00c9251",
  1607 => x"ab972d80",
  1608 => x"dc900880",
  1609 => x"2e8c3880",
  1610 => x"ddf00880",
  1611 => x"c00780dd",
  1612 => x"f00c9451",
  1613 => x"ab972d80",
  1614 => x"dc900880",
  1615 => x"2e8b3880",
  1616 => x"ddf00890",
  1617 => x"0780ddf0",
  1618 => x"0c9151ab",
  1619 => x"972d80dc",
  1620 => x"9008802e",
  1621 => x"8b3880dd",
  1622 => x"f008a007",
  1623 => x"80ddf00c",
  1624 => x"9d51ab97",
  1625 => x"2d80dc90",
  1626 => x"08802e8b",
  1627 => x"3880ddf0",
  1628 => x"08810780",
  1629 => x"ddf00c9b",
  1630 => x"51ab972d",
  1631 => x"80dc9008",
  1632 => x"802e8b38",
  1633 => x"80ddf008",
  1634 => x"820780dd",
  1635 => x"f00c9c51",
  1636 => x"ab972d80",
  1637 => x"dc900880",
  1638 => x"2e8b3880",
  1639 => x"ddf00884",
  1640 => x"0780ddf0",
  1641 => x"0ca351ab",
  1642 => x"972d80dc",
  1643 => x"9008802e",
  1644 => x"8b3880dd",
  1645 => x"f0088807",
  1646 => x"80ddf00c",
  1647 => x"81fd51ab",
  1648 => x"972d81fa",
  1649 => x"51ab972d",
  1650 => x"b9a00481",
  1651 => x"f551ab97",
  1652 => x"2d80dc90",
  1653 => x"08812a70",
  1654 => x"81065152",
  1655 => x"71802eb3",
  1656 => x"3880ddfc",
  1657 => x"08527180",
  1658 => x"2e8a38ff",
  1659 => x"1280ddfc",
  1660 => x"0cb49304",
  1661 => x"80ddf808",
  1662 => x"1080ddf8",
  1663 => x"08057084",
  1664 => x"29165152",
  1665 => x"88120880",
  1666 => x"2e8938ff",
  1667 => x"51881208",
  1668 => x"52712d81",
  1669 => x"f251ab97",
  1670 => x"2d80dc90",
  1671 => x"08812a70",
  1672 => x"81065152",
  1673 => x"71802eb4",
  1674 => x"3880ddf8",
  1675 => x"08ff1180",
  1676 => x"ddfc0856",
  1677 => x"53537372",
  1678 => x"258a3881",
  1679 => x"1480ddfc",
  1680 => x"0cb4dc04",
  1681 => x"72101370",
  1682 => x"84291651",
  1683 => x"52881208",
  1684 => x"802e8938",
  1685 => x"fe518812",
  1686 => x"0852712d",
  1687 => x"81fd51ab",
  1688 => x"972d80dc",
  1689 => x"9008812a",
  1690 => x"70810651",
  1691 => x"5271802e",
  1692 => x"b13880dd",
  1693 => x"fc08802e",
  1694 => x"8a38800b",
  1695 => x"80ddfc0c",
  1696 => x"b5a20480",
  1697 => x"ddf80810",
  1698 => x"80ddf808",
  1699 => x"05708429",
  1700 => x"16515288",
  1701 => x"1208802e",
  1702 => x"8938fd51",
  1703 => x"88120852",
  1704 => x"712d81fa",
  1705 => x"51ab972d",
  1706 => x"80dc9008",
  1707 => x"812a7081",
  1708 => x"06515271",
  1709 => x"802eb138",
  1710 => x"80ddf808",
  1711 => x"ff115452",
  1712 => x"80ddfc08",
  1713 => x"73258938",
  1714 => x"7280ddfc",
  1715 => x"0cb5e804",
  1716 => x"71101270",
  1717 => x"84291651",
  1718 => x"52881208",
  1719 => x"802e8938",
  1720 => x"fc518812",
  1721 => x"0852712d",
  1722 => x"80ddfc08",
  1723 => x"70535473",
  1724 => x"802e8a38",
  1725 => x"8c15ff15",
  1726 => x"5555b5ef",
  1727 => x"04820b80",
  1728 => x"dca40c71",
  1729 => x"8f0680dc",
  1730 => x"a00c81eb",
  1731 => x"51ab972d",
  1732 => x"80dc9008",
  1733 => x"812a7081",
  1734 => x"06515271",
  1735 => x"802ead38",
  1736 => x"7408852e",
  1737 => x"098106a4",
  1738 => x"38881580",
  1739 => x"f52dff05",
  1740 => x"52718816",
  1741 => x"81b72d71",
  1742 => x"982b5271",
  1743 => x"80258838",
  1744 => x"800b8816",
  1745 => x"81b72d74",
  1746 => x"51adfc2d",
  1747 => x"81f451ab",
  1748 => x"972d80dc",
  1749 => x"9008812a",
  1750 => x"70810651",
  1751 => x"5271802e",
  1752 => x"b3387408",
  1753 => x"852e0981",
  1754 => x"06aa3888",
  1755 => x"1580f52d",
  1756 => x"81055271",
  1757 => x"881681b7",
  1758 => x"2d7181ff",
  1759 => x"068b1680",
  1760 => x"f52d5452",
  1761 => x"72722787",
  1762 => x"38728816",
  1763 => x"81b72d74",
  1764 => x"51adfc2d",
  1765 => x"80da51ab",
  1766 => x"972d80dc",
  1767 => x"9008812a",
  1768 => x"70810651",
  1769 => x"5271802e",
  1770 => x"81ad3880",
  1771 => x"ddf40880",
  1772 => x"ddfc0855",
  1773 => x"5373802e",
  1774 => x"8a388c13",
  1775 => x"ff155553",
  1776 => x"b7b50472",
  1777 => x"08527182",
  1778 => x"2ea63871",
  1779 => x"82268938",
  1780 => x"71812eaa",
  1781 => x"38b8d704",
  1782 => x"71832eb4",
  1783 => x"3871842e",
  1784 => x"09810680",
  1785 => x"f2388813",
  1786 => x"0851afd2",
  1787 => x"2db8d704",
  1788 => x"80ddfc08",
  1789 => x"51881308",
  1790 => x"52712db8",
  1791 => x"d704810b",
  1792 => x"8814082b",
  1793 => x"80dacc08",
  1794 => x"3280dacc",
  1795 => x"0cb8ab04",
  1796 => x"881380f5",
  1797 => x"2d81058b",
  1798 => x"1480f52d",
  1799 => x"53547174",
  1800 => x"24833880",
  1801 => x"54738814",
  1802 => x"81b72dae",
  1803 => x"ac2db8d7",
  1804 => x"04750880",
  1805 => x"2ea43875",
  1806 => x"0851ab97",
  1807 => x"2d80dc90",
  1808 => x"08810652",
  1809 => x"71802e8c",
  1810 => x"3880ddfc",
  1811 => x"08518416",
  1812 => x"0852712d",
  1813 => x"88165675",
  1814 => x"d8388054",
  1815 => x"800b80dc",
  1816 => x"a40c738f",
  1817 => x"0680dca0",
  1818 => x"0ca05273",
  1819 => x"80ddfc08",
  1820 => x"2e098106",
  1821 => x"993880dd",
  1822 => x"f808ff05",
  1823 => x"74327009",
  1824 => x"81057072",
  1825 => x"079f2a91",
  1826 => x"71315151",
  1827 => x"53537151",
  1828 => x"83842d81",
  1829 => x"14548e74",
  1830 => x"25c23880",
  1831 => x"dad00852",
  1832 => x"7180dc90",
  1833 => x"0c029805",
  1834 => x"0d0402f4",
  1835 => x"050dd452",
  1836 => x"81ff720c",
  1837 => x"71085381",
  1838 => x"ff720c72",
  1839 => x"882b83fe",
  1840 => x"80067208",
  1841 => x"7081ff06",
  1842 => x"51525381",
  1843 => x"ff720c72",
  1844 => x"7107882b",
  1845 => x"72087081",
  1846 => x"ff065152",
  1847 => x"5381ff72",
  1848 => x"0c727107",
  1849 => x"882b7208",
  1850 => x"7081ff06",
  1851 => x"720780dc",
  1852 => x"900c5253",
  1853 => x"028c050d",
  1854 => x"0402f405",
  1855 => x"0d747671",
  1856 => x"81ff06d4",
  1857 => x"0c535380",
  1858 => x"de840885",
  1859 => x"3871892b",
  1860 => x"5271982a",
  1861 => x"d40c7190",
  1862 => x"2a7081ff",
  1863 => x"06d40c51",
  1864 => x"71882a70",
  1865 => x"81ff06d4",
  1866 => x"0c517181",
  1867 => x"ff06d40c",
  1868 => x"72902a70",
  1869 => x"81ff06d4",
  1870 => x"0c51d408",
  1871 => x"7081ff06",
  1872 => x"515182b8",
  1873 => x"bf527081",
  1874 => x"ff2e0981",
  1875 => x"06943881",
  1876 => x"ff0bd40c",
  1877 => x"d4087081",
  1878 => x"ff06ff14",
  1879 => x"54515171",
  1880 => x"e5387080",
  1881 => x"dc900c02",
  1882 => x"8c050d04",
  1883 => x"02fc050d",
  1884 => x"81c75181",
  1885 => x"ff0bd40c",
  1886 => x"ff115170",
  1887 => x"8025f438",
  1888 => x"0284050d",
  1889 => x"0402f405",
  1890 => x"0d81ff0b",
  1891 => x"d40c9353",
  1892 => x"805287fc",
  1893 => x"80c151b9",
  1894 => x"f92d80dc",
  1895 => x"90088b38",
  1896 => x"81ff0bd4",
  1897 => x"0c8153bb",
  1898 => x"b304baec",
  1899 => x"2dff1353",
  1900 => x"72de3872",
  1901 => x"80dc900c",
  1902 => x"028c050d",
  1903 => x"0402ec05",
  1904 => x"0d810b80",
  1905 => x"de840c84",
  1906 => x"54d00870",
  1907 => x"8f2a7081",
  1908 => x"06515153",
  1909 => x"72f33872",
  1910 => x"d00cbaec",
  1911 => x"2d80d6dc",
  1912 => x"5186a02d",
  1913 => x"d008708f",
  1914 => x"2a708106",
  1915 => x"51515372",
  1916 => x"f338810b",
  1917 => x"d00cb153",
  1918 => x"805284d4",
  1919 => x"80c051b9",
  1920 => x"f92d80dc",
  1921 => x"9008812e",
  1922 => x"93387282",
  1923 => x"2ebf38ff",
  1924 => x"135372e4",
  1925 => x"38ff1454",
  1926 => x"73ffae38",
  1927 => x"baec2d83",
  1928 => x"aa52849c",
  1929 => x"80c851b9",
  1930 => x"f92d80dc",
  1931 => x"9008812e",
  1932 => x"09810693",
  1933 => x"38b9aa2d",
  1934 => x"80dc9008",
  1935 => x"83ffff06",
  1936 => x"537283aa",
  1937 => x"2e9f38bb",
  1938 => x"852dbce0",
  1939 => x"0480d6e8",
  1940 => x"5186a02d",
  1941 => x"8053beb5",
  1942 => x"0480d780",
  1943 => x"5186a02d",
  1944 => x"8054be86",
  1945 => x"0481ff0b",
  1946 => x"d40cb154",
  1947 => x"baec2d8f",
  1948 => x"cf538052",
  1949 => x"87fc80f7",
  1950 => x"51b9f92d",
  1951 => x"80dc9008",
  1952 => x"5580dc90",
  1953 => x"08812e09",
  1954 => x"81069c38",
  1955 => x"81ff0bd4",
  1956 => x"0c820a52",
  1957 => x"849c80e9",
  1958 => x"51b9f92d",
  1959 => x"80dc9008",
  1960 => x"802e8d38",
  1961 => x"baec2dff",
  1962 => x"135372c6",
  1963 => x"38bdf904",
  1964 => x"81ff0bd4",
  1965 => x"0c80dc90",
  1966 => x"085287fc",
  1967 => x"80fa51b9",
  1968 => x"f92d80dc",
  1969 => x"9008b238",
  1970 => x"81ff0bd4",
  1971 => x"0cd40853",
  1972 => x"81ff0bd4",
  1973 => x"0c81ff0b",
  1974 => x"d40c81ff",
  1975 => x"0bd40c81",
  1976 => x"ff0bd40c",
  1977 => x"72862a70",
  1978 => x"81067656",
  1979 => x"51537296",
  1980 => x"3880dc90",
  1981 => x"0854be86",
  1982 => x"0473822e",
  1983 => x"fedb38ff",
  1984 => x"145473fe",
  1985 => x"e7387380",
  1986 => x"de840c73",
  1987 => x"8b388152",
  1988 => x"87fc80d0",
  1989 => x"51b9f92d",
  1990 => x"81ff0bd4",
  1991 => x"0cd00870",
  1992 => x"8f2a7081",
  1993 => x"06515153",
  1994 => x"72f33872",
  1995 => x"d00c81ff",
  1996 => x"0bd40c81",
  1997 => x"537280dc",
  1998 => x"900c0294",
  1999 => x"050d0402",
  2000 => x"e8050d78",
  2001 => x"55805681",
  2002 => x"ff0bd40c",
  2003 => x"d008708f",
  2004 => x"2a708106",
  2005 => x"51515372",
  2006 => x"f3388281",
  2007 => x"0bd00c81",
  2008 => x"ff0bd40c",
  2009 => x"775287fc",
  2010 => x"80d151b9",
  2011 => x"f92d80db",
  2012 => x"c6df5480",
  2013 => x"dc900880",
  2014 => x"2e8b3880",
  2015 => x"d7a05186",
  2016 => x"a02dbfd9",
  2017 => x"0481ff0b",
  2018 => x"d40cd408",
  2019 => x"7081ff06",
  2020 => x"51537281",
  2021 => x"fe2e0981",
  2022 => x"069e3880",
  2023 => x"ff53b9aa",
  2024 => x"2d80dc90",
  2025 => x"08757084",
  2026 => x"05570cff",
  2027 => x"13537280",
  2028 => x"25ec3881",
  2029 => x"56bfbe04",
  2030 => x"ff145473",
  2031 => x"c83881ff",
  2032 => x"0bd40c81",
  2033 => x"ff0bd40c",
  2034 => x"d008708f",
  2035 => x"2a708106",
  2036 => x"51515372",
  2037 => x"f33872d0",
  2038 => x"0c7580dc",
  2039 => x"900c0298",
  2040 => x"050d0402",
  2041 => x"e8050d77",
  2042 => x"797b5855",
  2043 => x"55805372",
  2044 => x"7625a438",
  2045 => x"74708105",
  2046 => x"5680f52d",
  2047 => x"74708105",
  2048 => x"5680f52d",
  2049 => x"52527171",
  2050 => x"2e873881",
  2051 => x"5180c099",
  2052 => x"04811353",
  2053 => x"bfef0480",
  2054 => x"517080dc",
  2055 => x"900c0298",
  2056 => x"050d0402",
  2057 => x"ec050d76",
  2058 => x"5574802e",
  2059 => x"80c4389a",
  2060 => x"1580e02d",
  2061 => x"5180ced1",
  2062 => x"2d80dc90",
  2063 => x"0880dc90",
  2064 => x"0880e4b8",
  2065 => x"0c80dc90",
  2066 => x"08545480",
  2067 => x"e4940880",
  2068 => x"2e9b3894",
  2069 => x"1580e02d",
  2070 => x"5180ced1",
  2071 => x"2d80dc90",
  2072 => x"08902b83",
  2073 => x"fff00a06",
  2074 => x"70750751",
  2075 => x"537280e4",
  2076 => x"b80c80e4",
  2077 => x"b8085372",
  2078 => x"802e9e38",
  2079 => x"80e48c08",
  2080 => x"fe147129",
  2081 => x"80e4a008",
  2082 => x"0580e4bc",
  2083 => x"0c70842b",
  2084 => x"80e4980c",
  2085 => x"5480c1c8",
  2086 => x"0480e4a4",
  2087 => x"0880e4b8",
  2088 => x"0c80e4a8",
  2089 => x"0880e4bc",
  2090 => x"0c80e494",
  2091 => x"08802e8c",
  2092 => x"3880e48c",
  2093 => x"08842b53",
  2094 => x"80c1c304",
  2095 => x"80e4ac08",
  2096 => x"842b5372",
  2097 => x"80e4980c",
  2098 => x"0294050d",
  2099 => x"0402d805",
  2100 => x"0d800b80",
  2101 => x"e4940c84",
  2102 => x"54bbbd2d",
  2103 => x"80dc9008",
  2104 => x"802e9838",
  2105 => x"80de8852",
  2106 => x"8051bebf",
  2107 => x"2d80dc90",
  2108 => x"08802e87",
  2109 => x"38fe5480",
  2110 => x"c28304ff",
  2111 => x"14547380",
  2112 => x"24d73873",
  2113 => x"8e3880d7",
  2114 => x"b05186a0",
  2115 => x"2d735580",
  2116 => x"c7e10480",
  2117 => x"56810b80",
  2118 => x"e4c00c88",
  2119 => x"5380d7c4",
  2120 => x"5280debe",
  2121 => x"51bfe32d",
  2122 => x"80dc9008",
  2123 => x"762e0981",
  2124 => x"06893880",
  2125 => x"dc900880",
  2126 => x"e4c00c88",
  2127 => x"5380d7d0",
  2128 => x"5280deda",
  2129 => x"51bfe32d",
  2130 => x"80dc9008",
  2131 => x"893880dc",
  2132 => x"900880e4",
  2133 => x"c00c80e4",
  2134 => x"c008802e",
  2135 => x"81843880",
  2136 => x"e1ce0b80",
  2137 => x"f52d80e1",
  2138 => x"cf0b80f5",
  2139 => x"2d71982b",
  2140 => x"71902b07",
  2141 => x"80e1d00b",
  2142 => x"80f52d70",
  2143 => x"882b7207",
  2144 => x"80e1d10b",
  2145 => x"80f52d71",
  2146 => x"0780e286",
  2147 => x"0b80f52d",
  2148 => x"80e2870b",
  2149 => x"80f52d71",
  2150 => x"882b0753",
  2151 => x"5f54525a",
  2152 => x"56575573",
  2153 => x"81abaa2e",
  2154 => x"09810690",
  2155 => x"38755180",
  2156 => x"cea02d80",
  2157 => x"dc900856",
  2158 => x"80c3cb04",
  2159 => x"7382d4d5",
  2160 => x"2e893880",
  2161 => x"d7dc5180",
  2162 => x"c4980480",
  2163 => x"de885275",
  2164 => x"51bebf2d",
  2165 => x"80dc9008",
  2166 => x"5580dc90",
  2167 => x"08802e84",
  2168 => x"80388853",
  2169 => x"80d7d052",
  2170 => x"80deda51",
  2171 => x"bfe32d80",
  2172 => x"dc90088b",
  2173 => x"38810b80",
  2174 => x"e4940c80",
  2175 => x"c49f0488",
  2176 => x"5380d7c4",
  2177 => x"5280debe",
  2178 => x"51bfe32d",
  2179 => x"80dc9008",
  2180 => x"802e8c38",
  2181 => x"80d7f051",
  2182 => x"86a02d80",
  2183 => x"c4fe0480",
  2184 => x"e2860b80",
  2185 => x"f52d5473",
  2186 => x"80d52e09",
  2187 => x"810680ce",
  2188 => x"3880e287",
  2189 => x"0b80f52d",
  2190 => x"547381aa",
  2191 => x"2e098106",
  2192 => x"bd38800b",
  2193 => x"80de880b",
  2194 => x"80f52d56",
  2195 => x"547481e9",
  2196 => x"2e833881",
  2197 => x"547481eb",
  2198 => x"2e8c3880",
  2199 => x"5573752e",
  2200 => x"09810682",
  2201 => x"fc3880de",
  2202 => x"930b80f5",
  2203 => x"2d55748e",
  2204 => x"3880de94",
  2205 => x"0b80f52d",
  2206 => x"5473822e",
  2207 => x"87388055",
  2208 => x"80c7e104",
  2209 => x"80de950b",
  2210 => x"80f52d70",
  2211 => x"80e48c0c",
  2212 => x"ff0580e4",
  2213 => x"900c80de",
  2214 => x"960b80f5",
  2215 => x"2d80de97",
  2216 => x"0b80f52d",
  2217 => x"58760577",
  2218 => x"82802905",
  2219 => x"7080e49c",
  2220 => x"0c80de98",
  2221 => x"0b80f52d",
  2222 => x"7080e4b0",
  2223 => x"0c80e494",
  2224 => x"08595758",
  2225 => x"76802e81",
  2226 => x"b8388853",
  2227 => x"80d7d052",
  2228 => x"80deda51",
  2229 => x"bfe32d80",
  2230 => x"dc900882",
  2231 => x"843880e4",
  2232 => x"8c087084",
  2233 => x"2b80e498",
  2234 => x"0c7080e4",
  2235 => x"ac0c80de",
  2236 => x"ad0b80f5",
  2237 => x"2d80deac",
  2238 => x"0b80f52d",
  2239 => x"71828029",
  2240 => x"0580deae",
  2241 => x"0b80f52d",
  2242 => x"70848080",
  2243 => x"291280de",
  2244 => x"af0b80f5",
  2245 => x"2d708180",
  2246 => x"0a291270",
  2247 => x"80e4b40c",
  2248 => x"80e4b008",
  2249 => x"712980e4",
  2250 => x"9c080570",
  2251 => x"80e4a00c",
  2252 => x"80deb50b",
  2253 => x"80f52d80",
  2254 => x"deb40b80",
  2255 => x"f52d7182",
  2256 => x"80290580",
  2257 => x"deb60b80",
  2258 => x"f52d7084",
  2259 => x"80802912",
  2260 => x"80deb70b",
  2261 => x"80f52d70",
  2262 => x"982b81f0",
  2263 => x"0a067205",
  2264 => x"7080e4a4",
  2265 => x"0cfe117e",
  2266 => x"29770580",
  2267 => x"e4a80c52",
  2268 => x"59524354",
  2269 => x"5e515259",
  2270 => x"525d5759",
  2271 => x"5780c7d9",
  2272 => x"0480de9a",
  2273 => x"0b80f52d",
  2274 => x"80de990b",
  2275 => x"80f52d71",
  2276 => x"82802905",
  2277 => x"7080e498",
  2278 => x"0c70a029",
  2279 => x"83ff0570",
  2280 => x"892a7080",
  2281 => x"e4ac0c80",
  2282 => x"de9f0b80",
  2283 => x"f52d80de",
  2284 => x"9e0b80f5",
  2285 => x"2d718280",
  2286 => x"29057080",
  2287 => x"e4b40c7b",
  2288 => x"71291e70",
  2289 => x"80e4a80c",
  2290 => x"7d80e4a4",
  2291 => x"0c730580",
  2292 => x"e4a00c55",
  2293 => x"5e515155",
  2294 => x"55805180",
  2295 => x"c0a32d81",
  2296 => x"557480dc",
  2297 => x"900c02a8",
  2298 => x"050d0402",
  2299 => x"ec050d76",
  2300 => x"70872c71",
  2301 => x"80ff0655",
  2302 => x"565480e4",
  2303 => x"94088a38",
  2304 => x"73882c74",
  2305 => x"81ff0654",
  2306 => x"5580de88",
  2307 => x"5280e49c",
  2308 => x"081551be",
  2309 => x"bf2d80dc",
  2310 => x"90085480",
  2311 => x"dc900880",
  2312 => x"2ebb3880",
  2313 => x"e4940880",
  2314 => x"2e9c3872",
  2315 => x"842980de",
  2316 => x"88057008",
  2317 => x"525380ce",
  2318 => x"a02d80dc",
  2319 => x"9008f00a",
  2320 => x"065380c8",
  2321 => x"db047210",
  2322 => x"80de8805",
  2323 => x"7080e02d",
  2324 => x"525380ce",
  2325 => x"d12d80dc",
  2326 => x"90085372",
  2327 => x"547380dc",
  2328 => x"900c0294",
  2329 => x"050d0402",
  2330 => x"e0050d79",
  2331 => x"70842c80",
  2332 => x"e4bc0805",
  2333 => x"718f0652",
  2334 => x"5553728a",
  2335 => x"3880de88",
  2336 => x"527351be",
  2337 => x"bf2d72a0",
  2338 => x"2980de88",
  2339 => x"05548074",
  2340 => x"80f52d56",
  2341 => x"5374732e",
  2342 => x"83388153",
  2343 => x"7481e52e",
  2344 => x"81f53881",
  2345 => x"70740654",
  2346 => x"5872802e",
  2347 => x"81e9388b",
  2348 => x"1480f52d",
  2349 => x"70832a79",
  2350 => x"06585676",
  2351 => x"9c3880da",
  2352 => x"d4085372",
  2353 => x"89387280",
  2354 => x"e2880b81",
  2355 => x"b72d7680",
  2356 => x"dad40c73",
  2357 => x"5380cb99",
  2358 => x"04758f2e",
  2359 => x"09810681",
  2360 => x"b638749f",
  2361 => x"068d2980",
  2362 => x"e1fb1151",
  2363 => x"53811480",
  2364 => x"f52d7370",
  2365 => x"81055581",
  2366 => x"b72d8314",
  2367 => x"80f52d73",
  2368 => x"70810555",
  2369 => x"81b72d85",
  2370 => x"1480f52d",
  2371 => x"73708105",
  2372 => x"5581b72d",
  2373 => x"871480f5",
  2374 => x"2d737081",
  2375 => x"055581b7",
  2376 => x"2d891480",
  2377 => x"f52d7370",
  2378 => x"81055581",
  2379 => x"b72d8e14",
  2380 => x"80f52d73",
  2381 => x"70810555",
  2382 => x"81b72d90",
  2383 => x"1480f52d",
  2384 => x"73708105",
  2385 => x"5581b72d",
  2386 => x"921480f5",
  2387 => x"2d737081",
  2388 => x"055581b7",
  2389 => x"2d941480",
  2390 => x"f52d7370",
  2391 => x"81055581",
  2392 => x"b72d9614",
  2393 => x"80f52d73",
  2394 => x"70810555",
  2395 => x"81b72d98",
  2396 => x"1480f52d",
  2397 => x"73708105",
  2398 => x"5581b72d",
  2399 => x"9c1480f5",
  2400 => x"2d737081",
  2401 => x"055581b7",
  2402 => x"2d9e1480",
  2403 => x"f52d7381",
  2404 => x"b72d7780",
  2405 => x"dad40c80",
  2406 => x"537280dc",
  2407 => x"900c02a0",
  2408 => x"050d0402",
  2409 => x"cc050d7e",
  2410 => x"605e5a80",
  2411 => x"0b80e4b8",
  2412 => x"0880e4bc",
  2413 => x"08595c56",
  2414 => x"805880e4",
  2415 => x"9808782e",
  2416 => x"81bc3877",
  2417 => x"8f06a017",
  2418 => x"57547391",
  2419 => x"3880de88",
  2420 => x"52765181",
  2421 => x"1757bebf",
  2422 => x"2d80de88",
  2423 => x"56807680",
  2424 => x"f52d5654",
  2425 => x"74742e83",
  2426 => x"38815474",
  2427 => x"81e52e81",
  2428 => x"81388170",
  2429 => x"7506555c",
  2430 => x"73802e80",
  2431 => x"f5388b16",
  2432 => x"80f52d98",
  2433 => x"06597880",
  2434 => x"e9388b53",
  2435 => x"7c527551",
  2436 => x"bfe32d80",
  2437 => x"dc900880",
  2438 => x"d9389c16",
  2439 => x"085180ce",
  2440 => x"a02d80dc",
  2441 => x"9008841b",
  2442 => x"0c9a1680",
  2443 => x"e02d5180",
  2444 => x"ced12d80",
  2445 => x"dc900880",
  2446 => x"dc900888",
  2447 => x"1c0c80dc",
  2448 => x"90085555",
  2449 => x"80e49408",
  2450 => x"802e9a38",
  2451 => x"941680e0",
  2452 => x"2d5180ce",
  2453 => x"d12d80dc",
  2454 => x"9008902b",
  2455 => x"83fff00a",
  2456 => x"06701651",
  2457 => x"5473881b",
  2458 => x"0c787a0c",
  2459 => x"7b5480cd",
  2460 => x"bc048118",
  2461 => x"5880e498",
  2462 => x"087826fe",
  2463 => x"c63880e4",
  2464 => x"9408802e",
  2465 => x"b5387a51",
  2466 => x"80c7eb2d",
  2467 => x"80dc9008",
  2468 => x"80dc9008",
  2469 => x"80ffffff",
  2470 => x"f806555b",
  2471 => x"7380ffff",
  2472 => x"fff82e96",
  2473 => x"3880dc90",
  2474 => x"08fe0580",
  2475 => x"e48c0829",
  2476 => x"80e4a008",
  2477 => x"055780cb",
  2478 => x"b8048054",
  2479 => x"7380dc90",
  2480 => x"0c02b405",
  2481 => x"0d0402f4",
  2482 => x"050d7470",
  2483 => x"08810571",
  2484 => x"0c700880",
  2485 => x"e4900806",
  2486 => x"53537190",
  2487 => x"38881308",
  2488 => x"5180c7eb",
  2489 => x"2d80dc90",
  2490 => x"0888140c",
  2491 => x"810b80dc",
  2492 => x"900c028c",
  2493 => x"050d0402",
  2494 => x"f0050d75",
  2495 => x"881108fe",
  2496 => x"0580e48c",
  2497 => x"082980e4",
  2498 => x"a0081172",
  2499 => x"0880e490",
  2500 => x"08060579",
  2501 => x"55535454",
  2502 => x"bebf2d02",
  2503 => x"90050d04",
  2504 => x"02f4050d",
  2505 => x"7470882a",
  2506 => x"83fe8006",
  2507 => x"7072982a",
  2508 => x"0772882b",
  2509 => x"87fc8080",
  2510 => x"0673982b",
  2511 => x"81f00a06",
  2512 => x"71730707",
  2513 => x"80dc900c",
  2514 => x"56515351",
  2515 => x"028c050d",
  2516 => x"0402f805",
  2517 => x"0d028e05",
  2518 => x"80f52d74",
  2519 => x"882b0770",
  2520 => x"83ffff06",
  2521 => x"80dc900c",
  2522 => x"51028805",
  2523 => x"0d0402f4",
  2524 => x"050d7476",
  2525 => x"78535452",
  2526 => x"80712597",
  2527 => x"38727081",
  2528 => x"055480f5",
  2529 => x"2d727081",
  2530 => x"055481b7",
  2531 => x"2dff1151",
  2532 => x"70eb3880",
  2533 => x"7281b72d",
  2534 => x"028c050d",
  2535 => x"0402e805",
  2536 => x"0d775680",
  2537 => x"70565473",
  2538 => x"7624b738",
  2539 => x"80e49808",
  2540 => x"742eaf38",
  2541 => x"735180c8",
  2542 => x"e72d80dc",
  2543 => x"900880dc",
  2544 => x"90080981",
  2545 => x"057080dc",
  2546 => x"9008079f",
  2547 => x"2a770581",
  2548 => x"17575753",
  2549 => x"53747624",
  2550 => x"893880e4",
  2551 => x"98087426",
  2552 => x"d3387280",
  2553 => x"dc900c02",
  2554 => x"98050d04",
  2555 => x"02f0050d",
  2556 => x"80dc8c08",
  2557 => x"165180cf",
  2558 => x"9d2d80dc",
  2559 => x"9008802e",
  2560 => x"a0388b53",
  2561 => x"80dc9008",
  2562 => x"5280e288",
  2563 => x"5180ceee",
  2564 => x"2d80e4c4",
  2565 => x"08547380",
  2566 => x"2e873880",
  2567 => x"e2885173",
  2568 => x"2d029005",
  2569 => x"0d0402dc",
  2570 => x"050d8070",
  2571 => x"5a557480",
  2572 => x"dc8c0825",
  2573 => x"b53880e4",
  2574 => x"9808752e",
  2575 => x"ad387851",
  2576 => x"80c8e72d",
  2577 => x"80dc9008",
  2578 => x"09810570",
  2579 => x"80dc9008",
  2580 => x"079f2a76",
  2581 => x"05811b5b",
  2582 => x"56547480",
  2583 => x"dc8c0825",
  2584 => x"893880e4",
  2585 => x"98087926",
  2586 => x"d5388055",
  2587 => x"7880e498",
  2588 => x"082781e4",
  2589 => x"38785180",
  2590 => x"c8e72d80",
  2591 => x"dc900880",
  2592 => x"2e81b438",
  2593 => x"80dc9008",
  2594 => x"8b0580f5",
  2595 => x"2d70842a",
  2596 => x"70810677",
  2597 => x"1078842b",
  2598 => x"80e2880b",
  2599 => x"80f52d5c",
  2600 => x"5c535155",
  2601 => x"5673802e",
  2602 => x"80ce3874",
  2603 => x"16822b80",
  2604 => x"d2fc0b80",
  2605 => x"dae0120c",
  2606 => x"54777531",
  2607 => x"1080e4c8",
  2608 => x"11555690",
  2609 => x"74708105",
  2610 => x"5681b72d",
  2611 => x"a07481b7",
  2612 => x"2d7681ff",
  2613 => x"06811658",
  2614 => x"5473802e",
  2615 => x"8b389c53",
  2616 => x"80e28852",
  2617 => x"80d1ef04",
  2618 => x"8b5380dc",
  2619 => x"90085280",
  2620 => x"e4ca1651",
  2621 => x"80d2ad04",
  2622 => x"7416822b",
  2623 => x"80cfec0b",
  2624 => x"80dae012",
  2625 => x"0c547681",
  2626 => x"ff068116",
  2627 => x"58547380",
  2628 => x"2e8b389c",
  2629 => x"5380e288",
  2630 => x"5280d2a4",
  2631 => x"048b5380",
  2632 => x"dc900852",
  2633 => x"77753110",
  2634 => x"80e4c805",
  2635 => x"51765580",
  2636 => x"ceee2d80",
  2637 => x"d2cc0474",
  2638 => x"90297531",
  2639 => x"701080e4",
  2640 => x"c8055154",
  2641 => x"80dc9008",
  2642 => x"7481b72d",
  2643 => x"81195974",
  2644 => x"8b24a438",
  2645 => x"80d0ec04",
  2646 => x"74902975",
  2647 => x"31701080",
  2648 => x"e4c8058c",
  2649 => x"77315751",
  2650 => x"54807481",
  2651 => x"b72d9e14",
  2652 => x"ff165654",
  2653 => x"74f33802",
  2654 => x"a4050d04",
  2655 => x"02fc050d",
  2656 => x"80dc8c08",
  2657 => x"135180cf",
  2658 => x"9d2d80dc",
  2659 => x"9008802e",
  2660 => x"8a3880dc",
  2661 => x"90085180",
  2662 => x"c0a32d80",
  2663 => x"0b80dc8c",
  2664 => x"0c80d0a6",
  2665 => x"2daeac2d",
  2666 => x"0284050d",
  2667 => x"0402fc05",
  2668 => x"0d725170",
  2669 => x"fd2eb238",
  2670 => x"70fd248b",
  2671 => x"3870fc2e",
  2672 => x"80d03880",
  2673 => x"d49c0470",
  2674 => x"fe2eb938",
  2675 => x"70ff2e09",
  2676 => x"810680c8",
  2677 => x"3880dc8c",
  2678 => x"08517080",
  2679 => x"2ebe38ff",
  2680 => x"1180dc8c",
  2681 => x"0c80d49c",
  2682 => x"0480dc8c",
  2683 => x"08f00570",
  2684 => x"80dc8c0c",
  2685 => x"51708025",
  2686 => x"a338800b",
  2687 => x"80dc8c0c",
  2688 => x"80d49c04",
  2689 => x"80dc8c08",
  2690 => x"810580dc",
  2691 => x"8c0c80d4",
  2692 => x"9c0480dc",
  2693 => x"8c089005",
  2694 => x"80dc8c0c",
  2695 => x"80d0a62d",
  2696 => x"aeac2d02",
  2697 => x"84050d04",
  2698 => x"02fc050d",
  2699 => x"800b80dc",
  2700 => x"8c0c80d0",
  2701 => x"a62dada8",
  2702 => x"2d80dc90",
  2703 => x"0880dbfc",
  2704 => x"0c80dad8",
  2705 => x"51afd22d",
  2706 => x"0284050d",
  2707 => x"047180e4",
  2708 => x"c40c0400",
  2709 => x"00ffffff",
  2710 => x"ff00ffff",
  2711 => x"ffff00ff",
  2712 => x"ffffff00",
  2713 => x"30313233",
  2714 => x"34353637",
  2715 => x"38394142",
  2716 => x"43444546",
  2717 => x"00000000",
  2718 => x"44656275",
  2719 => x"67000000",
  2720 => x"52657365",
  2721 => x"74000000",
  2722 => x"5363616e",
  2723 => x"6c696e65",
  2724 => x"73000000",
  2725 => x"50414c20",
  2726 => x"2f204e54",
  2727 => x"53430000",
  2728 => x"436f6c6f",
  2729 => x"72000000",
  2730 => x"44696666",
  2731 => x"6963756c",
  2732 => x"74792041",
  2733 => x"00000000",
  2734 => x"44696666",
  2735 => x"6963756c",
  2736 => x"74792042",
  2737 => x"00000000",
  2738 => x"2a537570",
  2739 => x"65726368",
  2740 => x"69702069",
  2741 => x"6e206361",
  2742 => x"72747269",
  2743 => x"64676500",
  2744 => x"2a42616e",
  2745 => x"6b204530",
  2746 => x"00000000",
  2747 => x"53656c65",
  2748 => x"63740000",
  2749 => x"53746172",
  2750 => x"74000000",
  2751 => x"4c6f6164",
  2752 => x"20524f4d",
  2753 => x"20100000",
  2754 => x"45786974",
  2755 => x"00000000",
  2756 => x"524f4d20",
  2757 => x"6c6f6164",
  2758 => x"696e6720",
  2759 => x"6661696c",
  2760 => x"65640000",
  2761 => x"4f4b0000",
  2762 => x"496e6974",
  2763 => x"69616c69",
  2764 => x"7a696e67",
  2765 => x"20534420",
  2766 => x"63617264",
  2767 => x"0a000000",
  2768 => x"436f6c6c",
  2769 => x"6563746f",
  2770 => x"72566973",
  2771 => x"696f6e00",
  2772 => x"16200000",
  2773 => x"14200000",
  2774 => x"15200000",
  2775 => x"53442069",
  2776 => x"6e69742e",
  2777 => x"2e2e0a00",
  2778 => x"53442063",
  2779 => x"61726420",
  2780 => x"72657365",
  2781 => x"74206661",
  2782 => x"696c6564",
  2783 => x"210a0000",
  2784 => x"53444843",
  2785 => x"20657272",
  2786 => x"6f72210a",
  2787 => x"00000000",
  2788 => x"57726974",
  2789 => x"65206661",
  2790 => x"696c6564",
  2791 => x"0a000000",
  2792 => x"52656164",
  2793 => x"20666169",
  2794 => x"6c65640a",
  2795 => x"00000000",
  2796 => x"43617264",
  2797 => x"20696e69",
  2798 => x"74206661",
  2799 => x"696c6564",
  2800 => x"0a000000",
  2801 => x"46415431",
  2802 => x"36202020",
  2803 => x"00000000",
  2804 => x"46415433",
  2805 => x"32202020",
  2806 => x"00000000",
  2807 => x"4e6f2070",
  2808 => x"61727469",
  2809 => x"74696f6e",
  2810 => x"20736967",
  2811 => x"0a000000",
  2812 => x"42616420",
  2813 => x"70617274",
  2814 => x"0a000000",
  2815 => x"4261636b",
  2816 => x"00000000",
  2817 => x"00000002",
  2818 => x"00002a64",
  2819 => x"00002e7c",
  2820 => x"00000002",
  2821 => x"00002e38",
  2822 => x"000012e6",
  2823 => x"00000002",
  2824 => x"00002a78",
  2825 => x"00001276",
  2826 => x"00000002",
  2827 => x"00002a80",
  2828 => x"0000035a",
  2829 => x"00000001",
  2830 => x"00002a88",
  2831 => x"00000000",
  2832 => x"00000001",
  2833 => x"00002a94",
  2834 => x"00000001",
  2835 => x"00000001",
  2836 => x"00002aa0",
  2837 => x"00000002",
  2838 => x"00000001",
  2839 => x"00002aa8",
  2840 => x"00000003",
  2841 => x"00000001",
  2842 => x"00002ab8",
  2843 => x"00000004",
  2844 => x"00000001",
  2845 => x"00002ac8",
  2846 => x"00000005",
  2847 => x"00000001",
  2848 => x"00002ae0",
  2849 => x"00000008",
  2850 => x"00000002",
  2851 => x"00002aec",
  2852 => x"0000036e",
  2853 => x"00000002",
  2854 => x"00002af4",
  2855 => x"00000a3f",
  2856 => x"00000002",
  2857 => x"00002afc",
  2858 => x"00002a28",
  2859 => x"00000002",
  2860 => x"00002b08",
  2861 => x"000016c5",
  2862 => x"00000000",
  2863 => x"00000000",
  2864 => x"00000000",
  2865 => x"00000004",
  2866 => x"00002b10",
  2867 => x"00002cc4",
  2868 => x"00000004",
  2869 => x"00002b24",
  2870 => x"00002c10",
  2871 => x"00000000",
  2872 => x"00000000",
  2873 => x"00000000",
  2874 => x"00000000",
  2875 => x"00000000",
  2876 => x"00000000",
  2877 => x"00000000",
  2878 => x"00000000",
  2879 => x"00000000",
  2880 => x"00000000",
  2881 => x"00000000",
  2882 => x"00000000",
  2883 => x"00000000",
  2884 => x"00000000",
  2885 => x"00000000",
  2886 => x"00000000",
  2887 => x"00000000",
  2888 => x"00000000",
  2889 => x"00000000",
  2890 => x"00000000",
  2891 => x"76f55a1c",
  2892 => x"f21c1c1c",
  2893 => x"1c1c1c1c",
  2894 => x"00000000",
  2895 => x"00000fff",
  2896 => x"00000fff",
  2897 => x"00000000",
  2898 => x"00000000",
  2899 => x"00000006",
  2900 => x"00000000",
  2901 => x"00000000",
  2902 => x"00000002",
  2903 => x"00003248",
  2904 => x"000027ec",
  2905 => x"00000002",
  2906 => x"00003266",
  2907 => x"000027ec",
  2908 => x"00000002",
  2909 => x"00003284",
  2910 => x"000027ec",
  2911 => x"00000002",
  2912 => x"000032a2",
  2913 => x"000027ec",
  2914 => x"00000002",
  2915 => x"000032c0",
  2916 => x"000027ec",
  2917 => x"00000002",
  2918 => x"000032de",
  2919 => x"000027ec",
  2920 => x"00000002",
  2921 => x"000032fc",
  2922 => x"000027ec",
  2923 => x"00000002",
  2924 => x"0000331a",
  2925 => x"000027ec",
  2926 => x"00000002",
  2927 => x"00003338",
  2928 => x"000027ec",
  2929 => x"00000002",
  2930 => x"00003356",
  2931 => x"000027ec",
  2932 => x"00000002",
  2933 => x"00003374",
  2934 => x"000027ec",
  2935 => x"00000002",
  2936 => x"00003392",
  2937 => x"000027ec",
  2938 => x"00000002",
  2939 => x"000033b0",
  2940 => x"000027ec",
  2941 => x"00000004",
  2942 => x"00002bfc",
  2943 => x"00000000",
  2944 => x"00000000",
  2945 => x"00000000",
  2946 => x"000029ad",
  2947 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

